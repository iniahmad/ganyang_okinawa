`include "top_arrhythmia.v"

module top_arrhythmia_tb;

    // Parameters
    parameter BITSIZE = 20;

    // Inputs
    reg clk;
    reg reset;
    reg [BITSIZE*10-1:0] x;
    reg [6:0] test_index;
    // reg valid;

    // Outputs
    wire [BITSIZE-1:0] y1;
    wire [BITSIZE-1:0] y2;
    wire [BITSIZE*2-1:0] y;
    wire done_flag;
    // wire [BITSIZE-1:0] y2;

    // Instantiate the Unit Under Test (UUT)
    top_arrhythmia #(BITSIZE) uut (
        .clk(clk),
        .reset(reset),
        .x(x),
        .y({y1,y2}),
        .done_flag_out(done_flag)
    );

/// for output ///
    localparam max_data = 201;
    integer i;
    integer sum;
    integer true;
    logic pred  [max_data-1:0];
    logic reall [max_data-1:0];

    function logic compare_sign_mag;
        input [BITSIZE-1:0] val_a;
        input [BITSIZE-1:0] val_b;  // Declare inputs as 16-bit
        logic sign_a;
        logic sign_b;
        logic [BITSIZE-2:0] mag_a;
        logic [BITSIZE-2:0] mag_b;

        begin
            // Extract sign and magnitude
            sign_a = val_a[BITSIZE-1];
            sign_b = val_b[BITSIZE-1];
            mag_a = val_a[BITSIZE-2:0];
            mag_b = val_b[BITSIZE-2:0];

            // Compare based on sign and magnitude
            if (sign_a != sign_b) begin
                // If signs differ, the negative number is smaller
                compare_sign_mag = (sign_a < sign_b);  // 1 if A > B
            end else begin
                // If signs are the same, compare magnitudes
                if (sign_a == 1'b1) begin
                    // Both negative: larger magnitude means smaller number
                    compare_sign_mag = (mag_a < mag_b);  // 1 if (-)A > (-)B
                end else begin
                    // Both positive: larger magnitude means larger number
                    compare_sign_mag = (mag_a > mag_b);  // 1 if A > B
                end
            end
        end
    endfunction
/// for output ///

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10 time units period
    end

    // Test sequence
    initial begin
        $dumpfile("top_arrhythmia_tb.vcd");
        $dumpvars(0, top_arrhythmia_tb);
        // Initialize Inputs
        reset = 1;
        x = 0;

        // Wait for global reset to finish
        #10;
        reset = 0;

// Testcase 0 True
test_index = 16'd0;
x = {
20'b00000100001011000011,
20'b00000001111111000101,
20'b00000110010111111100,
20'b00000100011001110010,
20'b00000100001101110100,
20'b00000001010011110011,
20'b00000001010100101110,
20'b00000101111010011110,
20'b00000011101101100101,
20'b00000010101111111000
};
#600;
reall[0] = 1;

pred [0] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 1 False
test_index = 16'd1;
x = {
20'b00000100011100011100,
20'b00000011101101000010,
20'b00000011010010010100,
20'b00000011011010111011,
20'b00000010101011100001,
20'b00000100100110110010,
20'b00000010101001110011,
20'b00000100001100000100,
20'b00000011100110001001,
20'b00000011011010111011
};
#600;
reall[1] = 0;

pred [1] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 2 False
test_index = 16'd2;
x = {
20'b00000101110110111000,
20'b00000110000011011101,
20'b00000101111110011011,
20'b00000101110100010111,
20'b00000101101011100011,
20'b00000101101010010011,
20'b00000101100001011111,
20'b00000101101110000100,
20'b00000101110011000110,
20'b00000110000010001100
};
#600;
reall[2] = 0;

pred [2] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 3 True
test_index = 16'd3;
x = {
20'b00000011010101000100,
20'b00000010110110010001,
20'b00000010111010010101,
20'b00000011001011010101,
20'b00000010110100101010,
20'b00000010111001100001,
20'b00000011000011001111,
20'b00000010001100111101,
20'b00000100010111011111,
20'b00000011010001110100
};
#600;
reall[3] = 1;

pred [3] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 4 True
test_index = 16'd4;
x = {
20'b00000011101110110010,
20'b00000110010111101010,
20'b00000010111010000101,
20'b00000101101111110111,
20'b00000011010110000011,
20'b00000011000010101100,
20'b00000011000010101100,
20'b00000100101110010000,
20'b00000100100101101001,
20'b00000100110101110010
};
#600;
reall[4] = 1;

pred [4] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 5 False
test_index = 16'd5;
x = {
20'b00000101100110100001,
20'b00000101010010011001,
20'b00000101010110001011,
20'b00000101111101001010,
20'b00000110000000111100,
20'b00000101011110111110,
20'b00000101100100000000,
20'b00000101100110100001,
20'b00000101101011100011,
20'b00000101010001001000
};
#600;
reall[5] = 0;

pred [5] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 6 True
test_index = 16'd6;
x = {
20'b00000100011000111100,
20'b00000010101111111010,
20'b00001000000000000000,
20'b00000101111011011001,
20'b00000101110011100001,
20'b00000011110000001111,
20'b00000111100101101111,
20'b00000101111011011001,
20'b00000101110111011101,
20'b00000011101101100111
};
#600;
reall[6] = 1;

pred [6] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 7 True
test_index = 16'd7;
x = {
20'b00000100010110100101,
20'b00000011110110010100,
20'b00000011001011010010,
20'b00000100100110101110,
20'b00000001110010000001,
20'b00000001110011000101,
20'b00000111010010110100,
20'b00000011010110000011,
20'b00000101101101101101,
20'b00000011100010111101
};
#600;
reall[7] = 1;

pred [7] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 8 False
test_index = 16'd8;
x = {
20'b00000110010001000111,
20'b00000110010001000111,
20'b00000101100001010010,
20'b00000101011111000111,
20'b00000101111100011101,
20'b00000110000000110100,
20'b00000101111000000111,
20'b00000101010110011010,
20'b00000101111110101001,
20'b00000110010011010010
};
#600;
reall[8] = 0;

pred [8] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 9 False
test_index = 16'd9;
x = {
20'b00000110000011111110,
20'b00000101111010011011,
20'b00000101110000111001,
20'b00000110001011111011,
20'b00000110000111001001,
20'b00000101111111001101,
20'b00000101110101101010,
20'b00000101111111001101,
20'b00000101111000110110,
20'b00000110000011111110
};
#600;
reall[9] = 0;

pred [9] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 10 True
test_index = 16'd10;
x = {
20'b00000001011111011100,
20'b00000010000110110111,
20'b00000001110110010001,
20'b00000001110001000101,
20'b00000001101000010001,
20'b00000010101000000100,
20'b00000001100111101111,
20'b00000010000110110111,
20'b00000001110100001100,
20'b00000001100101001001
};
#600;
reall[10] = 1;

pred [10] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 11 True
test_index = 16'd11;
x = {
20'b00000010111101100100,
20'b00000011000100110111,
20'b00000001000110011110,
20'b00000001000110011110,
20'b00000100010010101000,
20'b00000011010111011111,
20'b00000001010011011100,
20'b00000000110011110110,
20'b00000011100010110101,
20'b00000011110010001110
};
#600;
reall[11] = 1;

pred [11] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 12 False
test_index = 16'd12;
x = {
20'b00000101111111101000,
20'b00000101111110001001,
20'b00000101111011001101,
20'b00000101111100101011,
20'b00000110001011011011,
20'b00000101111011001101,
20'b00000110000001000110,
20'b00000101110110110001,
20'b00000101110101010011,
20'b00000101111011001101
};
#600;
reall[12] = 0;

pred [12] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 13 False
test_index = 16'd13;
x = {
20'b00000100111011101101,
20'b00000101000000111010,
20'b00000100111100110000,
20'b00000101000000111010,
20'b00000100111110110101,
20'b00000100111111110111,
20'b00000101001100010101,
20'b00000100011100100011,
20'b00000101011011111010,
20'b00000101001111011100
};
#600;
reall[13] = 0;

pred [13] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 14 True
test_index = 16'd14;
x = {
20'b00000011000000110111,
20'b00000101100000000000,
20'b00000010111100100010,
20'b00000101000110111010,
20'b00000011110011111001,
20'b00000011100000110111,
20'b00000011110101100111,
20'b00000100101101110101,
20'b00000100011001000101,
20'b00000100011100100010
};
#600;
reall[14] = 1;

pred [14] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 15 False
test_index = 16'd15;
x = {
20'b00000101101111010011,
20'b00000101101000111100,
20'b00000101101100000111,
20'b00000101100010100101,
20'b00000101110000111001,
20'b00000101110010011111,
20'b00000101101100000111,
20'b00000101100010100101,
20'b00000101101000111100,
20'b00000101101010100010
};
#600;
reall[15] = 0;

pred [15] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 16 True
test_index = 16'd16;
x = {
20'b00000110001101011001,
20'b00000100111010000010,
20'b00000100101111101000,
20'b00000100110100000101,
20'b00000100101110001000,
20'b00000100110001000111,
20'b00000011000111011100,
20'b00000110011001010011,
20'b00000100011010110010,
20'b00000101001010011010
};
#600;
reall[16] = 1;

pred [16] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 17 False
test_index = 16'd17;
x = {
20'b00000101110011011010,
20'b00000101111010010110,
20'b00000101101101010101,
20'b00000101011011000111,
20'b00000101011101101110,
20'b00000101101111111100,
20'b00000101110111110000,
20'b00000101100110011001,
20'b00000101010111101001,
20'b00000101011100110110
};
#600;
reall[17] = 0;

pred [17] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 18 False
test_index = 16'd18;
x = {
20'b00000010110010001110,
20'b00000011001100111101,
20'b00000010111111001100,
20'b00000010110110010001,
20'b00000010111100110000,
20'b00000011101011101111,
20'b00000011010111011111,
20'b00000100001101110001,
20'b00000010101110001011,
20'b00000010110100101010
};
#600;
reall[18] = 0;

pred [18] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 19 False
test_index = 16'd19;
x = {
20'b00000101100100000000,
20'b00000101100101010001,
20'b00000101110100010111,
20'b00000101111001011001,
20'b00000101111110011011,
20'b00000101101100110100,
20'b00000101100001011111,
20'b00000101100000001111,
20'b00000101100100000000,
20'b00000101101110000100
};
#600;
reall[19] = 0;

pred [19] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 20 False
test_index = 16'd20;
x = {
20'b00000100111000100001,
20'b00000100101111011000,
20'b00000100111011110110,
20'b00000100111100101011,
20'b00000100101011001110,
20'b00000100111011000000,
20'b00000100110100010111,
20'b00000111001101010011,
20'b00000011101100111000,
20'b00000101011011011011
};
#600;
reall[20] = 0;

pred [20] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 21 False
test_index = 16'd21;
x = {
20'b00000101100000001110,
20'b00000101011110010111,
20'b00000110011011000110,
20'b00000110110100010100,
20'b00000110100111001111,
20'b00000111001001110011,
20'b00000110110100010100,
20'b00000101110011110110,
20'b00000110010111010110,
20'b00000110010110011011
};
#600;
reall[21] = 0;

pred [21] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 22 False
test_index = 16'd22;
x = {
20'b00000011010100111001,
20'b00000011010010010100,
20'b00000100011011100101,
20'b00000011101010011100,
20'b00000011100101010001,
20'b00000100000100010011,
20'b00000100110000010001,
20'b00000101000100000110,
20'b00000011100011100011,
20'b00000011100101010001
};
#600;
reall[22] = 0;

pred [22] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 23 False
test_index = 16'd23;
x = {
20'b00000101111111001011,
20'b00000101111010001110,
20'b00000101011001001011,
20'b00000110010111111100,
20'b00000101101110101010,
20'b00000110001010101111,
20'b00000110011001100110,
20'b00000110010100101001,
20'b00000110000100001000,
20'b00000101111111001011
};
#600;
reall[23] = 0;

pred [23] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 24 False
test_index = 16'd24;
x = {
20'b00000110000101100010,
20'b00000110000010100101,
20'b00000110000010100101,
20'b00000110001110011000,
20'b00000110001001111101,
20'b00000110000101100010,
20'b00000110001000011110,
20'b00000110010100010010,
20'b00000110010001010101,
20'b00000101111110001001
};
#600;
reall[24] = 0;

pred [24] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 25 False
test_index = 16'd25;
x = {
20'b00000100100111000011,
20'b00000100011110010111,
20'b00000100000111001110,
20'b00000100001000101011,
20'b00000100001011100100,
20'b00000100000100010101,
20'b00000100001101000001,
20'b00000100001101000001,
20'b00000100100001010000,
20'b00000011101011110000
};
#600;
reall[25] = 0;

pred [25] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 26 False
test_index = 16'd26;
x = {
20'b00000100011011011110,
20'b00000100011111110100,
20'b00000100100100001010,
20'b00000100101011011000,
20'b00000100100100001010,
20'b00000100011011011110,
20'b00000100001111111010,
20'b00000100001010000111,
20'b00000100001011100100,
20'b00000100010100001111
};
#600;
reall[26] = 0;

pred [26] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 27 False
test_index = 16'd27;
x = {
20'b00000010101010001000,
20'b00000011110001011010,
20'b00000011000100110111,
20'b00000011111000101101,
20'b00000010101100100011,
20'b00000010101010001000,
20'b00000010100001001101,
20'b00000010101011101111,
20'b00000011001000111010,
20'b00000011011101111110
};
#600;
reall[27] = 0;

pred [27] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 28 True
test_index = 16'd28;
x = {
20'b00000101000010111110,
20'b00000100110101100101,
20'b00000100111000100011,
20'b00000100101100101001,
20'b00000100111000100011,
20'b00000100011010110010,
20'b00000101010011010110,
20'b00000100111110100000,
20'b00000011010100110101,
20'b00000110011001010011
};
#600;
reall[28] = 1;

pred [28] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 29 False
test_index = 16'd29;
x = {
20'b00000101111000110110,
20'b00000110000000110010,
20'b00000110000111001001,
20'b00000101111010011011,
20'b00000101110101101010,
20'b00000101111101100111,
20'b00000110001000101111,
20'b00000101111010011011,
20'b00000101101100000111,
20'b00000101110000111001
};
#600;
reall[29] = 0;

pred [29] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 30 True
test_index = 16'd30;
x = {
20'b00000110000110110111,
20'b00000010111000100011,
20'b00000010101011010011,
20'b00000011011001101010,
20'b00000011000101110010,
20'b00000100011010111110,
20'b00000100100011011111,
20'b00000101001000011001,
20'b00000011000100110110,
20'b00000111001100111001
};
#600;
reall[30] = 1;

pred [30] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 31 True
test_index = 16'd31;
x = {
20'b00000001100101001100,
20'b00000011001100000110,
20'b00000001110100110000,
20'b00000100010010001010,
20'b00000011111110010001,
20'b00000010001011001111,
20'b00000011011000001101,
20'b00000011110011111001,
20'b00000010100000000000,
20'b00000011001000101001
};
#600;
reall[31] = 1;

pred [31] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 32 False
test_index = 16'd32;
x = {
20'b00000100110101110111,
20'b00000101001110011111,
20'b00000101100000111101,
20'b00000101101100001111,
20'b00000101010110101100,
20'b00000101010110101100,
20'b00000101010111101110,
20'b00000101000111010011,
20'b00000100110001110000,
20'b00000101000101010000
};
#600;
reall[32] = 0;

pred [32] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 33 False
test_index = 16'd33;
x = {
20'b00000110100100001011,
20'b00000110100001000100,
20'b00000110100100001011,
20'b00000110101000110110,
20'b00000110110110110110,
20'b00000111000000001100,
20'b00000110111101000101,
20'b00000110110010001100,
20'b00000110111110101000,
20'b00000111000111111110
};
#600;
reall[33] = 0;

pred [33] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 34 False
test_index = 16'd34;
x = {
20'b00000101011001110001,
20'b00000101100111000111,
20'b00000110001101000101,
20'b00000101011110111010,
20'b00000101011110111010,
20'b00000101111101101100,
20'b00000110111011010000,
20'b00000101111000100011,
20'b00000101110010011001,
20'b00000110001011000001
};
#600;
reall[34] = 0;

pred [34] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 35 False
test_index = 16'd35;
x = {
20'b00000101110010011111,
20'b00000101111111001101,
20'b00000110000101100100,
20'b00000101111100000001,
20'b00000101110010011111,
20'b00000101110111010000,
20'b00000101111000110110,
20'b00000110000011111110,
20'b00000110001000101111,
20'b00000101110101101010
};
#600;
reall[35] = 0;

pred [35] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 36 True
test_index = 16'd36;
x = {
20'b00000100111010011011,
20'b00000001011101111101,
20'b00000010100001011011,
20'b00000101100111000000,
20'b00000100010000010000,
20'b00000101011101010111,
20'b00000100011111111011,
20'b00000100111100110101,
20'b00000100011100010011,
20'b00000101000000011100
};
#600;
reall[36] = 1;

pred [36] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 37 False
test_index = 16'd37;
x = {
20'b00000100111000011010,
20'b00000100011111110100,
20'b00000100011000100101,
20'b00000100000111001110,
20'b00000100000101110010,
20'b00000100001000101011,
20'b00000100010010110011,
20'b00000100011100111011,
20'b00000100100111000011,
20'b00000100110100000100
};
#600;
reall[37] = 0;

pred [37] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 38 True
test_index = 16'd38;
x = {
20'b00000010101100001111,
20'b00000010101111000101,
20'b00000110000100111101,
20'b00000010010101100001,
20'b00000101110100111000,
20'b00000010100110100100,
20'b00000101110011111011,
20'b00000010111111001011,
20'b00000101100010111001,
20'b00000010110001111011
};
#600;
reall[38] = 1;

pred [38] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 39 False
test_index = 16'd39;
x = {
20'b00000100110010101100,
20'b00000100110011111101,
20'b00000100101110111001,
20'b00000100101001110100,
20'b00000100101110111001,
20'b00000100111001000001,
20'b00000100101100010110,
20'b00000100101011000101,
20'b00000100101001110100,
20'b00000100110001011011
};
#600;
reall[39] = 0;

pred [39] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 40 False
test_index = 16'd40;
x = {
20'b00000110001111111100,
20'b00000110001001101110,
20'b00000110000001111100,
20'b00000110010100100111,
20'b00000110010011000100,
20'b00000110001111111100,
20'b00000110000110100111,
20'b00000110010011000100,
20'b00000110001110011001,
20'b00000110001111111100
};
#600;
reall[40] = 0;

pred [40] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 41 False
test_index = 16'd41;
x = {
20'b00000101101100001111,
20'b00000101111011101000,
20'b00000110000000110001,
20'b00000101111011101000,
20'b00000101011010110011,
20'b00000110010000001010,
20'b00000110100110101110,
20'b00000110000111111100,
20'b00000101000010001011,
20'b00000101000011001101
};
#600;
reall[41] = 0;

pred [41] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 42 False
test_index = 16'd42;
x = {
20'b00000101101101010001,
20'b00000110000011110110,
20'b00000110000111111100,
20'b00000101011100110110,
20'b00000100111000111100,
20'b00000101100101000100,
20'b00000110010010001101,
20'b00000110011101011111,
20'b00000101110100011101,
20'b00000101111100101010
};
#600;
reall[42] = 0;

pred [42] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 43 True
test_index = 16'd43;
x = {
20'b00000010111011011010,
20'b00000111001110101110,
20'b00000010111100011000,
20'b00000111001001111001,
20'b00000010111010011100,
20'b00000111010000101010,
20'b00000010111100011000,
20'b00000011100010000011,
20'b00000011100011000001,
20'b00000100111011111001
};
#600;
reall[43] = 1;

pred [43] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 44 False
test_index = 16'd44;
x = {
20'b00000101100011110001,
20'b00000101101011101001,
20'b00000101101100111101,
20'b00000101100110011001,
20'b00000101101001000001,
20'b00000101101110010001,
20'b00000101100011110001,
20'b00000101101001000001,
20'b00000101011110100001,
20'b00000101011101001101
};
#600;
reall[44] = 0;

pred [44] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 45 False
test_index = 16'd45;
x = {
20'b00000111010000100011,
20'b00000111001000110100,
20'b00000111011001011000,
20'b00000111010111001011,
20'b00000111001011000010,
20'b00000111011101110010,
20'b00000111001011000010,
20'b00000111010010110000,
20'b00000111000111101110,
20'b00000111010000100011
};
#600;
reall[45] = 0;

pred [45] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 46 False
test_index = 16'd46;
x = {
20'b00000110000001111010,
20'b00000110000101101110,
20'b00000110010111100011,
20'b00000110101010101010,
20'b00000110101001011001,
20'b00000110010001001100,
20'b00000110000111000000,
20'b00000110010110010010,
20'b00000110100110110110,
20'b00000110100110110110
};
#600;
reall[46] = 0;

pred [46] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 47 True
test_index = 16'd47;
x = {
20'b00000111110101100101,
20'b00000110010011001010,
20'b00000010110010110111,
20'b00000010100001110101,
20'b00000111011010001001,
20'b00000110011001110010,
20'b00000011000001000100,
20'b00000010101101001100,
20'b00000111101001010010,
20'b00000110001001101100
};
#600;
reall[47] = 1;

pred [47] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 48 False
test_index = 16'd48;
x = {
20'b00000100110101001001,
20'b00000100111010000001,
20'b00000100110011001100,
20'b00000100101100010111,
20'b00000100110001001111,
20'b00000100110111000110,
20'b00000100101001011100,
20'b00000100100110100001,
20'b00000100101111010011,
20'b00000100101001011100
};
#600;
reall[48] = 0;

pred [48] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 49 False
test_index = 16'd49;
x = {
20'b00000011010101011110,
20'b00000011000100000111,
20'b00000010100000100010,
20'b00000011110101100101,
20'b00000011111001111011,
20'b00000100000110000100,
20'b00000010011001100110,
20'b00000100000110111100,
20'b00000010001111001011,
20'b00000100010100110100
};
#600;
reall[49] = 0;

pred [49] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 50 True
test_index = 16'd50;
x = {
20'b00000111000110111111,
20'b00000011111000011110,
20'b00000101110010000001,
20'b00000011101011100100,
20'b00000100100011011111,
20'b00000011000001100111,
20'b00000101011000001100,
20'b00000011101000010101,
20'b00000100111011001010,
20'b00000011100111010000
};
#600;
reall[50] = 1;

pred [50] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 51 True
test_index = 16'd51;
x = {
20'b00000001101111100100,
20'b00000011010101100111,
20'b00000011011011101011,
20'b00000011011001000101,
20'b00000010000000110111,
20'b00000101110011000001,
20'b00000010000001101110,
20'b00000011101101110101,
20'b00000011011001111100,
20'b00000011000000000000
};
#600;
reall[51] = 1;

pred [51] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 52 False
test_index = 16'd52;
x = {
20'b00000110010111100011,
20'b00000110000101101110,
20'b00000110001100000110,
20'b00000110001000010001,
20'b00000110100001110000,
20'b00000110011101111011,
20'b00000110101010101010,
20'b00000110100101100100,
20'b00000110000101101110,
20'b00000110001101010111
};
#600;
reall[52] = 0;

pred [52] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 53 True
test_index = 16'd53;
x = {
20'b00000011110000111100,
20'b00000100001100111010,
20'b00000001101000010101,
20'b00000001101000010101,
20'b00000100011001110100,
20'b00000011001101011100,
20'b00000100110010100011,
20'b00000011001101011100,
20'b00000100110010100011,
20'b00000011011101100101
};
#600;
reall[53] = 1;

pred [53] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 54 False
test_index = 16'd54;
x = {
20'b00000010100011001001,
20'b00000011110101100101,
20'b00000011011111000001,
20'b00000101000111001010,
20'b00000010110000001010,
20'b00000010110000001010,
20'b00000010101010111101,
20'b00000010111011011100,
20'b00000011101110101001,
20'b00000010111110111010
};
#600;
reall[54] = 0;

pred [54] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 55 False
test_index = 16'd55;
x = {
20'b00000100100100101111,
20'b00000100111011101000,
20'b00000100100100101111,
20'b00000100100100101111,
20'b00000100100001001000,
20'b00000100101001100011,
20'b00000100100101111100,
20'b00000100101001100011,
20'b00000100100100101111,
20'b00000100100100101111
};
#600;
reall[55] = 0;

pred [55] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 56 False
test_index = 16'd56;
x = {
20'b00000101110101101010,
20'b00000101101111010011,
20'b00000101101100000111,
20'b00000101100100001011,
20'b00000101101010100010,
20'b00000101100111010110,
20'b00000101110010011111,
20'b00000101111000110110,
20'b00000101100111010110,
20'b00000101100100001011
};
#600;
reall[56] = 0;

pred [56] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 57 False
test_index = 16'd57;
x = {
20'b00000100100110000001,
20'b00000100101011000101,
20'b00000100100111010010,
20'b00000100110001011011,
20'b00000100110010101100,
20'b00000100101101100111,
20'b00000100100010001101,
20'b00000100100111010010,
20'b00000100101101100111,
20'b00000100101101100111
};
#600;
reall[57] = 0;

pred [57] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 58 False
test_index = 16'd58;
x = {
20'b00000101110111010000,
20'b00000101111010011011,
20'b00000110000000110010,
20'b00000110000011111110,
20'b00000110000011111110,
20'b00000101111100000001,
20'b00000101111000110110,
20'b00000101111101100111,
20'b00000110001011111011,
20'b00000110000000110010
};
#600;
reall[58] = 0;

pred [58] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 59 False
test_index = 16'd59;
x = {
20'b00000101110010101011,
20'b00000110101001000010,
20'b00000101101110010101,
20'b00000101100011011101,
20'b00000110001100110001,
20'b00000110000010111111,
20'b00000101011001101011,
20'b00000101000011111100,
20'b00000101110001100110,
20'b00000101101101001111
};
#600;
reall[59] = 0;

pred [59] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 60 True
test_index = 16'd60;
x = {
20'b00000001110101100111,
20'b00000001101100111110,
20'b00000011101001100000,
20'b00000010000101001100,
20'b00000010100111110010,
20'b00000010111101011001,
20'b00000010111011101011,
20'b00000011010110011111,
20'b00000010001111100100,
20'b00000010001000101001
};
#600;
reall[60] = 1;

pred [60] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 61 True
test_index = 16'd61;
x = {
20'b00000100000111101001,
20'b00000010000100101011,
20'b00000100010101010000,
20'b00000010000001010001,
20'b00000100010000001010,
20'b00000001111011000010,
20'b00000100010000001010,
20'b00000010000110111100,
20'b00000100010101110101,
20'b00000001111111000000
};
#600;
reall[61] = 1;

pred [61] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 62 False
test_index = 16'd62;
x = {
20'b00000101001111111001,
20'b00000101011000100110,
20'b00000101100010011000,
20'b00000101011010110001,
20'b00000101110010101011,
20'b00000111000110011000,
20'b00000110011011111111,
20'b00000110010101011110,
20'b00000110000010111111,
20'b00000101110001100110
};
#600;
reall[62] = 0;

pred [62] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 63 False
test_index = 16'd63;
x = {
20'b00000011001110110111,
20'b00000011110011000100,
20'b00000100010000011000,
20'b00000100010000011000,
20'b00000100001110101001,
20'b00000100011100011100,
20'b00000011010110101000,
20'b00000011101101000010,
20'b00000011001000110101,
20'b00000011111111001000
};
#600;
reall[63] = 0;

pred [63] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 64 False
test_index = 16'd64;
x = {
20'b00000101101010010011,
20'b00000101101001000010,
20'b00000101100000001111,
20'b00000101111110011011,
20'b00000110000111001110,
20'b00000101011101101110,
20'b00000101010100111010,
20'b00000101100110100001,
20'b00000101110001110110,
20'b00000101110000100101
};
#600;
reall[64] = 0;

pred [64] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 65 False
test_index = 16'd65;
x = {
20'b00000101110000010011,
20'b00000101110000010011,
20'b00000101100100101111,
20'b00000101110110111010,
20'b00000110001110000010,
20'b00000110010010111111,
20'b00000110000000110100,
20'b00000101110110111010,
20'b00000101111000100100,
20'b00000101111011110111
};
#600;
reall[65] = 0;

pred [65] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 66 False
test_index = 16'd66;
x = {
20'b00000110000001000110,
20'b00000101111000010000,
20'b00000110001001111101,
20'b00000101111100101011,
20'b00000110000101100010,
20'b00000110001100111010,
20'b00000110000101100010,
20'b00000110000101100010,
20'b00000110001111110111,
20'b00000110001011011011
};
#600;
reall[66] = 0;

pred [66] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 67 False
test_index = 16'd67;
x = {
20'b00000100100100011011,
20'b00000100111110111011,
20'b00000101000110100000,
20'b00000100110011100101,
20'b00000100100011011111,
20'b00000100100111010001,
20'b00000100101110110110,
20'b00000101000000110100,
20'b00000101010100101100,
20'b00000101010100101100
};
#600;
reall[67] = 0;

pred [67] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 68 False
test_index = 16'd68;
x = {
20'b00000110010100010000,
20'b00000101110011011011,
20'b00000101010001100100,
20'b00000110010101010010,
20'b00000110001000111110,
20'b00000101100111000111,
20'b00000110000110111011,
20'b00000101111111101111,
20'b00000110010010001101,
20'b00000101101100001111
};
#600;
reall[68] = 0;

pred [68] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 69 False
test_index = 16'd69;
x = {
20'b00000110001010111000,
20'b00000110000101010011,
20'b00000110011110111101,
20'b00000110100011011010,
20'b00000110011001011000,
20'b00000110010010101011,
20'b00000110001010111000,
20'b00000110001000101001,
20'b00000110010011110011,
20'b00000110110100001001
};
#600;
reall[69] = 0;

pred [69] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 70 True
test_index = 16'd70;
x = {
20'b00000001111001011000,
20'b00000001110100101101,
20'b00000001011110011010,
20'b00000010000110110111,
20'b00000001100111101111,
20'b00000001101100011010,
20'b00000001101111100001,
20'b00000001101101111110,
20'b00000010000100110011,
20'b00000001110011101011
};
#600;
reall[70] = 1;

pred [70] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 71 False
test_index = 16'd71;
x = {
20'b00000100001010111001,
20'b00000010100100000101,
20'b00000010011101110110,
20'b00000010110000100011,
20'b00000010101011010110,
20'b00000010010111101000,
20'b00000011101000101000,
20'b00000010111000110111,
20'b00000011000001001010,
20'b00000011011111010010
};
#600;
reall[71] = 0;

pred [71] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 72 False
test_index = 16'd72;
x = {
20'b00000100001011100100,
20'b00000100100001010000,
20'b00000100011000100101,
20'b00000100101011011000,
20'b00000100100101100110,
20'b00000100100101100110,
20'b00000100000111001110,
20'b00000100001011100100,
20'b00000100000010111001,
20'b00000100001101000001
};
#600;
reall[72] = 0;

pred [72] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 73 False
test_index = 16'd73;
x = {
20'b00000110011101011011,
20'b00000110100001100010,
20'b00000110111010001011,
20'b00000110111010001011,
20'b00000110111000110100,
20'b00000110010101001110,
20'b00000110000110001010,
20'b00000101111101111100,
20'b00000110001101000000,
20'b00000110101101110111
};
#600;
reall[73] = 0;

pred [73] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 74 False
test_index = 16'd74;
x = {
20'b00000101101100000111,
20'b00000101110100000100,
20'b00000101101111010011,
20'b00000101111100000001,
20'b00000101110111010000,
20'b00000101110111010000,
20'b00000101101010100010,
20'b00000101111111001101,
20'b00000101111010011011,
20'b00000101110101101010
};
#600;
reall[74] = 0;

pred [74] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 75 False
test_index = 16'd75;
x = {
20'b00000110110000110011,
20'b00000110110101010000,
20'b00000110010011110011,
20'b00000110011011100110,
20'b00000110010100111010,
20'b00000110010110000001,
20'b00000110100010010011,
20'b00000110110100001001,
20'b00000110101010000110,
20'b00000110001011111111
};
#600;
reall[75] = 0;

pred [75] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 76 False
test_index = 16'd76;
x = {
20'b00000110010011000100,
20'b00000110100001000100,
20'b00000110010111101110,
20'b00000110011010110110,
20'b00000110011111100000,
20'b00000110101010011010,
20'b00000110011001010010,
20'b00000110011100011001,
20'b00000110011111100000,
20'b00000110011111100000
};
#600;
reall[76] = 0;

pred [76] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 77 False
test_index = 16'd77;
x = {
20'b00000100110101001000,
20'b00000100110011001100,
20'b00000100110110000110,
20'b00000100111000111111,
20'b00000100110001010001,
20'b00000100101101011001,
20'b00000100111001111101,
20'b00000100111000111111,
20'b00000100110000010011,
20'b00000100111001111101
};
#600;
reall[77] = 0;

pred [77] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 78 False
test_index = 16'd78;
x = {
20'b00000100100111001001,
20'b00000100101000010110,
20'b00000100110001111111,
20'b00000100101010110001,
20'b00000100100011100010,
20'b00000100011110101110,
20'b00000100101001100011,
20'b00000100101001100011,
20'b00000100101010110001,
20'b00000011010000011010
};
#600;
reall[78] = 0;

pred [78] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 79 True
test_index = 16'd79;
x = {
20'b00000001101001010011,
20'b00000010000111011001,
20'b00000001110100001100,
20'b00000001101010010101,
20'b00000001001010001011,
20'b00000001001010001011,
20'b00000001110101001111,
20'b00000001011110011010,
20'b00000001011011110100,
20'b00000010011101101100
};
#600;
reall[79] = 1;

pred [79] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 80 False
test_index = 16'd80;
x = {
20'b00000101001111111001,
20'b00000101101000111001,
20'b00000101111101100011,
20'b00000101001111111001,
20'b00000100111110100000,
20'b00000101001100101000,
20'b00000101001110110011,
20'b00000101001100101000,
20'b00000100111100010101,
20'b00000101000010110110
};
#600;
reall[80] = 0;

pred [80] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 81 False
test_index = 16'd81;
x = {
20'b00000101100100000000,
20'b00000101100110100001,
20'b00000101101011100011,
20'b00000101010001001000,
20'b00000101011100011101,
20'b00000101101010010011,
20'b00000101110101100111,
20'b00000101100010110000,
20'b00000101010100111010,
20'b00000101000010000010
};
#600;
reall[81] = 0;

pred [81] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 82 False
test_index = 16'd82;
x = {
20'b00000101100111000111,
20'b00000101101110010011,
20'b00000101101101010001,
20'b00000101011000110000,
20'b00000101001111100001,
20'b00000100100110011110,
20'b00000100011100001101,
20'b00000100100100011011,
20'b00000101110101011110,
20'b00000110000001110010
};
#600;
reall[82] = 0;

pred [82] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 83 False
test_index = 16'd83;
x = {
20'b00000110000011100000,
20'b00000110000110100111,
20'b00000110000110100111,
20'b00000110000011100000,
20'b00000110000000011000,
20'b00000101111101010001,
20'b00000110001100110101,
20'b00000110000110100111,
20'b00000110000101000011,
20'b00000101111000100110
};
#600;
reall[83] = 0;

pred [83] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 84 False
test_index = 16'd84;
x = {
20'b00000110101011001110,
20'b00000110100001001011,
20'b00000110010001100100,
20'b00000101111010001001,
20'b00000101111100010111,
20'b00000101111110100110,
20'b00000110000110011010,
20'b00000101101110111111,
20'b00000101110110110011,
20'b00000101111011010000
};
#600;
reall[84] = 0;

pred [84] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 85 True
test_index = 16'd85;
x = {
20'b00000110011100111111,
20'b00000110010100100000,
20'b00000101001111001101,
20'b00000110111001010010,
20'b00000111000011001011,
20'b00000111000110000000,
20'b00000110110000110010,
20'b00000110011011100101,
20'b00000100111001111111,
20'b00000110101001101110
};
#600;
reall[85] = 1;

pred [85] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 86 False
test_index = 16'd86;
x = {
20'b00000100011010101111,
20'b00000100100010011000,
20'b00000100001100010011,
20'b00000100010010010000,
20'b00000100010000100011,
20'b00000100000010111110,
20'b00000100010011000110,
20'b00000100100001100010,
20'b00000100011111110101,
20'b00000100000010000111
};
#600;
reall[86] = 0;

pred [86] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 87 False
test_index = 16'd87;
x = {
20'b00000101101010100010,
20'b00000101110111010000,
20'b00000101110000111001,
20'b00000101111000110110,
20'b00000101111000110110,
20'b00000101110000111001,
20'b00000101100111010110,
20'b00000101111000110110,
20'b00000101111101100111,
20'b00000101110111010000
};
#600;
reall[87] = 0;

pred [87] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 88 True
test_index = 16'd88;
x = {
20'b00000100111010000010,
20'b00000001101001101011,
20'b00000001101001101011,
20'b00000110010000010111,
20'b00000100010011010110,
20'b00000101010111110100,
20'b00000011110100000101,
20'b00000011000000000000,
20'b00000011000001011111,
20'b00000100111000100011
};
#600;
reall[88] = 1;

pred [88] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 89 False
test_index = 16'd89;
x = {
20'b00000101100111101000,
20'b00000101101010011110,
20'b00000101001111000001,
20'b00000101100011110110,
20'b00000101011111000111,
20'b00000101101100010111,
20'b00000101000101100011,
20'b00000101010000111010,
20'b00000101111111010010,
20'b00000101110000001001
};
#600;
reall[89] = 0;

pred [89] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 90 False
test_index = 16'd90;
x = {
20'b00000101110111010000,
20'b00000101111010011011,
20'b00000101110010011111,
20'b00000101100101110000,
20'b00000101101101101101,
20'b00000101101101101101,
20'b00000101110010011111,
20'b00000101110101101010,
20'b00000101101000111100,
20'b00000101101000111100
};
#600;
reall[90] = 0;

pred [90] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 91 False
test_index = 16'd91;
x = {
20'b00000001011011100000,
20'b00000010010000101101,
20'b00000001011110011110,
20'b00000000111001011101,
20'b00000001101010011001,
20'b00000001010110011001,
20'b00000010000100010111,
20'b00000010010101110011,
20'b00000010010010110101,
20'b00000010001100011100
};
#600;
reall[91] = 0;

pred [91] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 92 False
test_index = 16'd92;
x = {
20'b00000101101100011100,
20'b00000101110000111000,
20'b00000101101100011100,
20'b00000101110000111000,
20'b00000101101001011111,
20'b00000101101000000001,
20'b00000101110010010110,
20'b00000101110011110100,
20'b00000101101000000001,
20'b00000101100011100110
};
#600;
reall[92] = 0;

pred [92] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 93 False
test_index = 16'd93;
x = {
20'b00000100110101001110,
20'b00000100111001000001,
20'b00000100110010101100,
20'b00000100101100010110,
20'b00000100110011111101,
20'b00000100111111010111,
20'b00000100110010101100,
20'b00000100110000001010,
20'b00000100110000001010,
20'b00000100110011111101
};
#600;
reall[93] = 0;

pred [93] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 94 False
test_index = 16'd94;
x = {
20'b00000111011110111001,
20'b00000111101100001000,
20'b00000111010010110000,
20'b00000111100111101110,
20'b00000111011100101100,
20'b00000111101110010110,
20'b00000111100000000000,
20'b00000111011110111001,
20'b00000111011011100101,
20'b00000111001110010110
};
#600;
reall[94] = 0;

pred [94] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 95 True
test_index = 16'd95;
x = {
20'b00000110110101001111,
20'b00000010100111100000,
20'b00000110100010010011,
20'b00000010101000011101,
20'b00000010011100001001,
20'b00000110111010111010,
20'b00000001011110101000,
20'b00000001011110101000,
20'b00000110111001111101,
20'b00000010101001011001
};
#600;
reall[95] = 1;

pred [95] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 96 False
test_index = 16'd96;
x = {
20'b00000101101100011100,
20'b00000101110110110001,
20'b00000101111100101011,
20'b00000101111011001101,
20'b00000101101010111110,
20'b00000110000001000110,
20'b00000101110010010110,
20'b00000101110110110001,
20'b00000101111111101000,
20'b00000101111011001101
};
#600;
reall[96] = 0;

pred [96] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 97 True
test_index = 16'd97;
x = {
20'b00000110110101100111,
20'b00000100101111010101,
20'b00000010111100011000,
20'b00000110101111110100,
20'b00000100110000010011,
20'b00000001101011001110,
20'b00000001100001100100,
20'b00000110100111000111,
20'b00000010110101100111,
20'b00000111001110101110
};
#600;
reall[97] = 1;

pred [97] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 98 False
test_index = 16'd98;
x = {
20'b00000100011101100000,
20'b00000100011000101100,
20'b00000100101111100101,
20'b00000100010111011111,
20'b00000100010101000101,
20'b00000100010011111000,
20'b00000100100111001001,
20'b00000100011110101110,
20'b00000100100011100010,
20'b00000100011101100000
};
#600;
reall[98] = 0;

pred [98] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 99 False
test_index = 16'd99;
x = {
20'b00000101001001100000,
20'b00000101001100000010,
20'b00000101001000001111,
20'b00000101000101101100,
20'b00000101000101101100,
20'b00000101001110100100,
20'b00000101001000001111,
20'b00000100111111010111,
20'b00000101000000101000,
20'b00000101001000001111
};
#600;
reall[99] = 0;

pred [99] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 100 False
test_index = 16'd100;
x = {
20'b00000101101110000100,
20'b00000101100110100001,
20'b00000101011101101110,
20'b00000101011110111110,
20'b00000101101010010011,
20'b00000101111010101001,
20'b00000101111000001000,
20'b00000101100110100001,
20'b00000101100110100001,
20'b00000101011011001101
};
#600;
reall[100] = 0;

pred [100] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 101 False
test_index = 16'd101;
x = {
20'b00000100010001101000,
20'b00000100010000011010,
20'b00000100100000001110,
20'b00000100011010001001,
20'b00000100100000001110,
20'b00000100101001111101,
20'b00000100101110110100,
20'b00000100100110010011,
20'b00000100011111000000,
20'b00000100010000011010
};
#600;
reall[101] = 0;

pred [101] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 102 False
test_index = 16'd102;
x = {
20'b00000010011001101101,
20'b00000100010010001011,
20'b00000010111010111011,
20'b00000011001010100000,
20'b00000100110001010101,
20'b00000100111011101101,
20'b00000011001100100101,
20'b00000010110011101010,
20'b00000100111000100110,
20'b00000010101001010010
};
#600;
reall[102] = 0;

pred [102] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 103 False
test_index = 16'd103;
x = {
20'b00000101111100000001,
20'b00000101110000111001,
20'b00000101111000110110,
20'b00000101110101101010,
20'b00000101111100000001,
20'b00000110000111001001,
20'b00000101111010011011,
20'b00000101110010011111,
20'b00000101111111001101,
20'b00000110001011111011
};
#600;
reall[103] = 0;

pred [103] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 104 False
test_index = 16'd104;
x = {
20'b00000101100011111101,
20'b00000101011110000111,
20'b00000101011010001101,
20'b00000101010110010011,
20'b00000101100000000011,
20'b00000101101000110101,
20'b00000101100000000011,
20'b00000101011011001011,
20'b00000101100110111000,
20'b00000101100101111010
};
#600;
reall[104] = 0;

pred [104] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 105 False
test_index = 16'd105;
x = {
20'b00000101011011110101,
20'b00000101011000110000,
20'b00000110100011101001,
20'b00000110010110010100,
20'b00000101011001110001,
20'b00000101010000100010,
20'b00000101001110011111,
20'b00000101011010110011,
20'b00000101100011000000,
20'b00000101011111111011
};
#600;
reall[105] = 0;

pred [105] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 106 False
test_index = 16'd106;
x = {
20'b00000110000001100101,
20'b00000110001001001010,
20'b00000110001100111101,
20'b00000110001010011011,
20'b00000110001110001110,
20'b00000110000111111001,
20'b00000110001110001110,
20'b00000101111011010000,
20'b00000101111001111111,
20'b00000110010011010001
};
#600;
reall[106] = 0;

pred [106] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 107 False
test_index = 16'd107;
x = {
20'b00000001110010111010,
20'b00000001100110100100,
20'b00000001010100101100,
20'b00000001010111101011,
20'b00000001011110111010,
20'b00000001100100011100,
20'b00000001001011110000,
20'b00000001010010001001,
20'b00000001001010011110,
20'b00000001100101010010
};
#600;
reall[107] = 0;

pred [107] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 108 False
test_index = 16'd108;
x = {
20'b00000101111000100011,
20'b00000110010100010000,
20'b00000110010011001111,
20'b00000101111101101100,
20'b00000101101010001100,
20'b00000101110011011011,
20'b00000110010100010000,
20'b00000101110011011011,
20'b00000101010001100100,
20'b00000110010101010010
};
#600;
reall[108] = 0;

pred [108] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 109 False
test_index = 16'd109;
x = {
20'b00000101101010110010,
20'b00000101100100111011,
20'b00000101100000000011,
20'b00000101011111000101,
20'b00000101011101001000,
20'b00000101100101111010,
20'b00000101100010111111,
20'b00000101100000000011,
20'b00000101100010111111,
20'b00000101100001000010
};
#600;
reall[109] = 0;

pred [109] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 110 False
test_index = 16'd110;
x = {
20'b00000100100110111100,
20'b00000100111001101000,
20'b00000100100111111110,
20'b00000100010100010000,
20'b00000101000001111100,
20'b00000100010100010000,
20'b00000100110011011010,
20'b00000100110010010111,
20'b00000100101111010000,
20'b00000100101101001011
};
#600;
reall[110] = 0;

pred [110] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 111 True
test_index = 16'd111;
x = {
20'b00000100011100111011,
20'b00000011001010011111,
20'b00000101101000001000,
20'b00000100001010000111,
20'b00000100001010000111,
20'b00000100000010111001,
20'b00000100000010111001,
20'b00000010100001111111,
20'b00000101111010111100,
20'b00000100011000100101
};
#600;
reall[111] = 1;

pred [111] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 112 True
test_index = 16'd112;
x = {
20'b00000010011001001101,
20'b00000011010111010110,
20'b00000010111110001111,
20'b00000010010001111110,
20'b00000001100010101111,
20'b00000001100010101111,
20'b00000010110011100110,
20'b00000001010101111110,
20'b00000011011110100101,
20'b00000010110100000001
};
#600;
reall[112] = 1;

pred [112] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 113 True
test_index = 16'd113;
x = {
20'b00000100001000010010,
20'b00000100000010110000,
20'b00000100000111010111,
20'b00000010100011111010,
20'b00000010101110111101,
20'b00001000000000000000,
20'b00000100010111000001,
20'b00000010100110101011,
20'b00000101010110100011,
20'b00000100000110011100
};
#600;
reall[113] = 1;

pred [113] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 114 False
test_index = 16'd114;
x = {
20'b00000110001010111000,
20'b00000110000111100001,
20'b00000110010110000001,
20'b00000110001011111111,
20'b00000101110100100100,
20'b00000110000100001011,
20'b00000110000101010011,
20'b00000101111110100110,
20'b00000110001010111000,
20'b00000101111111101110
};
#600;
reall[114] = 0;

pred [114] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 115 True
test_index = 16'd115;
x = {
20'b00000100110111000100,
20'b00000011010001110111,
20'b00000110010100110101,
20'b00000011111000100011,
20'b00000101111110100000,
20'b00000100111110100000,
20'b00000100110111000100,
20'b00000100110010100110,
20'b00000100110111000100,
20'b00000011011111010000
};
#600;
reall[115] = 1;

pred [115] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 116 True
test_index = 16'd116;
x = {
20'b00000110000011111010,
20'b00000011011110110111,
20'b00000110001000101110,
20'b00000011011011010000,
20'b00000101111001000100,
20'b00000011011101101010,
20'b00000110000110010100,
20'b00000011100111010011,
20'b00000101111101111001,
20'b00000011010010110100
};
#600;
reall[116] = 1;

pred [116] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 117 False
test_index = 16'd117;
x = {
20'b00000100011100010000,
20'b00000100011011011011,
20'b00000100100100100100,
20'b00000100100010111010,
20'b00000100010000100111,
20'b00000100001110001000,
20'b00000100001001111110,
20'b00000100011001110001,
20'b00000100010110011100,
20'b00000100011010100110
};
#600;
reall[117] = 0;

pred [117] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 118 False
test_index = 16'd118;
x = {
20'b00000111000010010101,
20'b00000101101011011100,
20'b00000101010001010010,
20'b00000101010010001110,
20'b00000101001101100011,
20'b00000101011110010111,
20'b00000101110011110110,
20'b00000111001100100111,
20'b00000111010011001001,
20'b00000111010111110100
};
#600;
reall[118] = 0;

pred [118] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 119 False
test_index = 16'd119;
x = {
20'b00000110001110011001,
20'b00000110000000011000,
20'b00000110000011100000,
20'b00000110000011100000,
20'b00000110001011010010,
20'b00000110000001111100,
20'b00000110000001111100,
20'b00000110000011100000,
20'b00000110001111111100,
20'b00000101111110110101
};
#600;
reall[119] = 0;

pred [119] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 120 False
test_index = 16'd120;
x = {
20'b00000101111010010110,
20'b00000101101101010101,
20'b00000101011011000111,
20'b00000101011101101110,
20'b00000101101111111100,
20'b00000101110111110000,
20'b00000101100110011001,
20'b00000101010111101001,
20'b00000101011100110110,
20'b00000101110110000001
};
#600;
reall[120] = 0;

pred [120] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 121 True
test_index = 16'd121;
x = {
20'b00000010011111010000,
20'b00000001110101110000,
20'b00000001010111101010,
20'b00000010111011110010,
20'b00000001100110001100,
20'b00000010010000001101,
20'b00000001110011101011,
20'b00000001110001000101,
20'b00000001010111001001,
20'b00000010001110101001
};
#600;
reall[121] = 1;

pred [121] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 122 True
test_index = 16'd122;
x = {
20'b00000011001010010110,
20'b00000100011010000011,
20'b00000010111011000001,
20'b00000101000100111110,
20'b00000010100011100000,
20'b00000011010111101000,
20'b00000101001100001000,
20'b00000010101000100111,
20'b00000001111011101010,
20'b00000100111101110101
};
#600;
reall[122] = 1;

pred [122] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 123 False
test_index = 16'd123;
x = {
20'b00000110011011100110,
20'b00000110010001100100,
20'b00000110011001011000,
20'b00000110010111001001,
20'b00000101111110100110,
20'b00000110000001111100,
20'b00000110101000111111,
20'b00000110100111111000,
20'b00000110001110001110,
20'b00000110001000101001
};
#600;
reall[123] = 0;

pred [123] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 124 False
test_index = 16'd124;
x = {
20'b00000111011110111001,
20'b00000111010111001011,
20'b00000111100001000110,
20'b00000111011000010001,
20'b00000111011110111001,
20'b00000111001100001000,
20'b00000111011001011000,
20'b00000111011100101100,
20'b00000111001001111011,
20'b00000111000110100111
};
#600;
reall[124] = 0;

pred [124] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 125 False
test_index = 16'd125;
x = {
20'b00000110001010110100,
20'b00000101111011100010,
20'b00000110001000010001,
20'b00000101110111101110,
20'b00000101110001010110,
20'b00000110001100000110,
20'b00000110011101111011,
20'b00000110001101010111,
20'b00000101110101001011,
20'b00000110000101101110
};
#600;
reall[125] = 0;

pred [125] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 126 False
test_index = 16'd126;
x = {
20'b00000100001000101011,
20'b00000100000010111001,
20'b00000100010001010110,
20'b00000100100100001010,
20'b00000100100100001010,
20'b00000100110010100111,
20'b00000100100100001010,
20'b00000100101001111100,
20'b00000100011011011110,
20'b00000100011011011110
};
#600;
reall[126] = 0;

pred [126] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 127 True
test_index = 16'd127;
x = {
20'b00000100001000101001,
20'b00000010100010100110,
20'b00000101001110101100,
20'b00000100000000000000,
20'b00000010011001000101,
20'b00000110001000101001,
20'b00000100100000000000,
20'b00000011111011101011,
20'b00000011110011000001,
20'b00000011111110010001
};
#600;
reall[127] = 1;

pred [127] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 128 False
test_index = 16'd128;
x = {
20'b00000011110111000101,
20'b00000011110001111111,
20'b00000011110001111111,
20'b00000100000010111110,
20'b00000011111011010101,
20'b00000100000010000111,
20'b00000011111011010101,
20'b00000011111000110010,
20'b00000011110110001111,
20'b00000011110110001111
};
#600;
reall[128] = 0;

pred [128] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 129 False
test_index = 16'd129;
x = {
20'b00000100010110011010,
20'b00000100000000000000,
20'b00000100011011100101,
20'b00000100000010100101,
20'b00000011110101101010,
20'b00000100010010111101,
20'b00000011110101101010,
20'b00000011111001111101,
20'b00000100001110101001,
20'b00000011110101101010
};
#600;
reall[129] = 0;

pred [129] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 130 False
test_index = 16'd130;
x = {
20'b00000011111010011000,
20'b00000100000111101010,
20'b00000011100001110110,
20'b00000011100001110110,
20'b00000011110010001101,
20'b00000100011110001001,
20'b00000011111010011000,
20'b00000100010000110111,
20'b00000011101101000110,
20'b00000011100010110111
};
#600;
reall[130] = 0;

pred [130] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 131 True
test_index = 16'd131;
x = {
20'b00000001001110110110,
20'b00000010110100000000,
20'b00000001100110101101,
20'b00000010011100001001,
20'b00000001110010000111,
20'b00000001010101000100,
20'b00000010101100001110,
20'b00000001100110001100,
20'b00000010100011011001,
20'b00000001111011011101
};
#600;
reall[131] = 1;

pred [131] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 132 False
test_index = 16'd132;
x = {
20'b00000011010110101000,
20'b00000010100111001110,
20'b00000011100101010001,
20'b00000010100011110001,
20'b00000010111010001011,
20'b00000011100111000000,
20'b00000011010100111001,
20'b00000011011000010110,
20'b00000011110110100001,
20'b00000011000111111110
};
#600;
reall[132] = 0;

pred [132] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 133 False
test_index = 16'd133;
x = {
20'b00000101110011011010,
20'b00000101101010101111,
20'b00000101010001100100,
20'b00000101011101101110,
20'b00000101101111111100,
20'b00000101111101110101,
20'b00000101101011100110,
20'b00000101011011111111,
20'b00000101101011100110,
20'b00000101110010100011
};
#600;
reall[133] = 0;

pred [133] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 134 False
test_index = 16'd134;
x = {
20'b00000110001100111010,
20'b00000110000100000011,
20'b00000110000010100101,
20'b00000101111110001001,
20'b00000110000010100101,
20'b00000101111110001001,
20'b00000110000101100010,
20'b00000110000101100010,
20'b00000101111110001001,
20'b00000101111000010000
};
#600;
reall[134] = 0;

pred [134] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 135 False
test_index = 16'd135;
x = {
20'b00000101011100011101,
20'b00000101011110111110,
20'b00000110000010001100,
20'b00000101110110111000,
20'b00000101110011000110,
20'b00000101101001000010,
20'b00000101100010110000,
20'b00000101100100000000,
20'b00000101101100110100,
20'b00000101100111110010
};
#600;
reall[135] = 0;

pred [135] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 136 True
test_index = 16'd136;
x = {
20'b00000100100111110011,
20'b00000100100011011111,
20'b00000011111011101100,
20'b00000011111101110110,
20'b00000100000000000000,
20'b00000001100101000110,
20'b00000001100101000110,
20'b00000100011011111101,
20'b00000011001111100110,
20'b00000101000100110101
};
#600;
reall[136] = 1;

pred [136] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 137 False
test_index = 16'd137;
x = {
20'b00000101111110100110,
20'b00000101111011010000,
20'b00000110010000011101,
20'b00000110101010000110,
20'b00000110100000000100,
20'b00000110010111001001,
20'b00000110011001011000,
20'b00000110010011110011,
20'b00000110001111010101,
20'b00000110101110100100
};
#600;
reall[137] = 0;

pred [137] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 138 False
test_index = 16'd138;
x = {
20'b00000101001011010010,
20'b00000101000111001011,
20'b00000101001000100011,
20'b00000101010010001000,
20'b00000101001011010010,
20'b00000101010011100000,
20'b00000101010000110001,
20'b00000101011111110101,
20'b00000101100010100100,
20'b00000011010100001100
};
#600;
reall[138] = 0;

pred [138] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 139 True
test_index = 16'd139;
x = {
20'b00000100010111000001,
20'b00000100000000111010,
20'b00000100000101100001,
20'b00000010000000111010,
20'b00000110010010011010,
20'b00000100100010000100,
20'b00000100100010111111,
20'b00000010010110000110,
20'b00000110000001110101,
20'b00000011110110110010
};
#600;
reall[139] = 1;

pred [139] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 140 True
test_index = 16'd140;
x = {
20'b00000101111101111000,
20'b00000110000011100010,
20'b00000110110011100111,
20'b00000100011100010010,
20'b00000110111110111100,
20'b00000111000000010110,
20'b00000110000010000111,
20'b00000100100110001100,
20'b00000111000111011011,
20'b00000110000110010111
};
#600;
reall[140] = 1;

pred [140] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 141 False
test_index = 16'd141;
x = {
20'b00000110010100111010,
20'b00000110000001111100,
20'b00000101110000000110,
20'b00000110000001111100,
20'b00000101101100110000,
20'b00000101101101110111,
20'b00000101101010100001,
20'b00000110000011000100,
20'b00000110100011011010,
20'b00000110001000101001
};
#600;
reall[141] = 0;

pred [141] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 142 True
test_index = 16'd142;
x = {
20'b00000011100110001101,
20'b00000011100110001101,
20'b00000010010111000001,
20'b00000100111101101100,
20'b00000011101101100101,
20'b00000011111000101000,
20'b00000011111001100011,
20'b00000011110100000001,
20'b00000010100000001110,
20'b00000100011111010011
};
#600;
reall[142] = 1;

pred [142] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 143 False
test_index = 16'd143;
x = {
20'b00000110001101000110,
20'b00000110001000101001,
20'b00000110000101010011,
20'b00000110000111100001,
20'b00000101110000000110,
20'b00000101111100010111,
20'b00000101110001001110,
20'b00000101100110000100,
20'b00000110001010111000,
20'b00000110100011011010
};
#600;
reall[143] = 0;

pred [143] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 144 True
test_index = 16'd144;
x = {
20'b00000100101000011010,
20'b00000101100001011111,
20'b00000100111110100111,
20'b00000100111101000001,
20'b00000101001100111000,
20'b00000101010011001110,
20'b00000100111011011100,
20'b00000101000110100010,
20'b00000101000001110010,
20'b00000100111001110110
};
#600;
reall[144] = 1;

pred [144] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 145 True
test_index = 16'd145;
x = {
20'b00000110001110111000,
20'b00000011011100010001,
20'b00000101110101100101,
20'b00000101000000000000,
20'b00000100111011100010,
20'b00000101000001011111,
20'b00000100110111000100,
20'b00000100110100000101,
20'b00000100111010000010,
20'b00000101000000000000
};
#600;
reall[145] = 1;

pred [145] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 146 False
test_index = 16'd146;
x = {
20'b00000101001110001000,
20'b00000101001110001000,
20'b00000100111100101011,
20'b00000101000110101001,
20'b00000100110101001100,
20'b00000101010010010010,
20'b00000101001101010011,
20'b00000100110111101100,
20'b00000100110101001100,
20'b00000100111000100001
};
#600;
reall[146] = 0;

pred [146] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 147 False
test_index = 16'd147;
x = {
20'b00000100100001100111,
20'b00000010101001110011,
20'b00000100100101111011,
20'b00000010110000101100,
20'b00000011110000011111,
20'b00000011100001110101,
20'b00000010100110010110,
20'b00000011010111011111,
20'b00000010111111010110,
20'b00000100001100111011
};
#600;
reall[147] = 0;

pred [147] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 148 True
test_index = 16'd148;
x = {
20'b00000110000111100001,
20'b00000011010100000001,
20'b00000110000101000111,
20'b00000011010100000001,
20'b00000101111010010001,
20'b00000011011000110110,
20'b00000110000101000111,
20'b00000011010111101001,
20'b00000101111011011110,
20'b00000011010100000001
};
#600;
reall[148] = 1;

pred [148] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 149 True
test_index = 16'd149;
x = {
20'b00000011010001001110,
20'b00000001010101100111,
20'b00000000111000001000,
20'b00000001011001100101,
20'b00000001001110001111,
20'b00000001010101100111,
20'b00000000111101001111,
20'b00000001010001000101,
20'b00000000001101100110,
20'b00000001110100001111
};
#600;
reall[149] = 1;

pred [149] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 150 False
test_index = 16'd150;
x = {
20'b00000100101110111001,
20'b00000100110101001110,
20'b00000100101110111001,
20'b00000100110110011111,
20'b00000100111100110101,
20'b00000100110011111101,
20'b00000100101110111001,
20'b00000100110101001110,
20'b00000100111010010011,
20'b00000100110111110000
};
#600;
reall[150] = 0;

pred [150] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 151 False
test_index = 16'd151;
x = {
20'b00000110000001111010,
20'b00000101111100110100,
20'b00000101111011100010,
20'b00000101101110110011,
20'b00000101101000011100,
20'b00000101110011111001,
20'b00000110001000010001,
20'b00000110001110101001,
20'b00000101111111010111,
20'b00000101111110000101
};
#600;
reall[151] = 0;

pred [151] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 152 False
test_index = 16'd152;
x = {
20'b00000011011001101011,
20'b00000011011011101110,
20'b00000100010101111110,
20'b00000011110101010001,
20'b00000110011000110010,
20'b00000100001010101110,
20'b00000100010000110111,
20'b00000100000111101010,
20'b00000011001101011010,
20'b00000011110111010100
};
#600;
reall[152] = 0;

pred [152] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 153 True
test_index = 16'd153;
x = {
20'b00000010001100001001,
20'b00000100000101101010,
20'b00000010111011001000,
20'b00000011101001010100,
20'b00000011001110100101,
20'b00000010101111110011,
20'b00000011001011010101,
20'b00000011110110010001,
20'b00000010000000110011,
20'b00000100101110111111
};
#600;
reall[153] = 1;

pred [153] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 154 True
test_index = 16'd154;
x = {
20'b00000000111110010001,
20'b00000010011100100010,
20'b00000010111000001101,
20'b00000100000001101110,
20'b00000100010011111001,
20'b00000001111001111100,
20'b00000001110001010011,
20'b00000011100000110111,
20'b00000011111010110011,
20'b00000100011101011001
};
#600;
reall[154] = 1;

pred [154] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 155 False
test_index = 16'd155;
x = {
20'b00000100101000101111,
20'b00000100101100011000,
20'b00000100101000101111,
20'b00000100100010101010,
20'b00000100101011001011,
20'b00000100111100001100,
20'b00000100111110101000,
20'b00000100111000100011,
20'b00000100101001111101,
20'b00000100101001111101
};
#600;
reall[155] = 0;

pred [155] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 156 True
test_index = 16'd156;
x = {
20'b00000100110001000111,
20'b00000100110100000101,
20'b00000011010110010100,
20'b00000110010110010100,
20'b00000101000101111101,
20'b00000100110111000100,
20'b00000011011010110010,
20'b00000110010001110111,
20'b00000101000100011101,
20'b00000100111110100000
};
#600;
reall[156] = 1;

pred [156] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 157 False
test_index = 16'd157;
x = {
20'b00000100011101001001,
20'b00000100011010100111,
20'b00000100011001010110,
20'b00000100010110110011,
20'b00000100011011111000,
20'b00000100011010100111,
20'b00000100010110110011,
20'b00000100010101100010,
20'b00000100010011000000,
20'b00000100011011111000
};
#600;
reall[157] = 0;

pred [157] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 158 False
test_index = 16'd158;
x = {
20'b00000110011010001010,
20'b00000110111000111111,
20'b00000111001011101011,
20'b00000110111101101010,
20'b00000111000111111100,
20'b00000101100110110001,
20'b00000101100111101101,
20'b00000101100111101101,
20'b00000101011011100011,
20'b00000101110000000111
};
#600;
reall[158] = 0;

pred [158] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 159 False
test_index = 16'd159;
x = {
20'b00000101000110111110,
20'b00000101001001100000,
20'b00000101001010110001,
20'b00000101001101010011,
20'b00000101001000001111,
20'b00000101000101101100,
20'b00000101000100011011,
20'b00000101010100111010,
20'b00000101001101010011,
20'b00000101000101101100
};
#600;
reall[159] = 0;

pred [159] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 160 False
test_index = 16'd160;
x = {
20'b00000110011001011000,
20'b00000110011110111101,
20'b00000110011101110101,
20'b00000110011010011111,
20'b00000110100101101001,
20'b00000110010100111010,
20'b00000101111011010000,
20'b00000101101100110000,
20'b00000101111110100110,
20'b00000110010100111010
};
#600;
reall[160] = 0;

pred [160] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 161 False
test_index = 16'd161;
x = {
20'b00000110110010110000,
20'b00000110111010011110,
20'b00000110110110000100,
20'b00000111000110100111,
20'b00000111001111011100,
20'b00000111011011100101,
20'b00000111010100111101,
20'b00000111100100011010,
20'b00000111011100101100,
20'b00000111011101110010
};
#600;
reall[161] = 0;

pred [161] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 162 True
test_index = 16'd162;
x = {
20'b00000010010110011011,
20'b00000001111000110111,
20'b00000001100111001110,
20'b00000010010010010010,
20'b00000001111110100100,
20'b00000001100101001001,
20'b00000010001011000001,
20'b00000001111000110111,
20'b00000001101100111011,
20'b00000010010111111111
};
#600;
reall[162] = 1;

pred [162] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 163 False
test_index = 16'd163;
x = {
20'b00000100101100000011,
20'b00000100011000000110,
20'b00000100011000111011,
20'b00000100110110110110,
20'b00000101010001011101,
20'b00000100011010100110,
20'b00000100111110010101,
20'b00000100110011100010,
20'b00000100011100010000,
20'b00000101001100011101
};
#600;
reall[163] = 0;

pred [163] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 164 True
test_index = 16'd164;
x = {
20'b00000100110001111011,
20'b00000100101110110000,
20'b00000100110011100001,
20'b00000100111000010001,
20'b00000100101011100101,
20'b00000100111101000001,
20'b00000100111011011100,
20'b00000100111001110110,
20'b00000100101110110000,
20'b00000100111011011100
};
#600;
reall[164] = 1;

pred [164] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 165 False
test_index = 16'd165;
x = {
20'b00000101111111010100,
20'b00000101110100010111,
20'b00000101011011101110,
20'b00000101001111011001,
20'b00000101010110001111,
20'b00000101101000000010,
20'b00000101111000011110,
20'b00000110000111100001,
20'b00000110000111100001,
20'b00000110001010010001
};
#600;
reall[165] = 0;

pred [165] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 166 False
test_index = 16'd166;
x = {
20'b00000110010000001010,
20'b00000110001100000011,
20'b00000101011000110000,
20'b00000101001111100001,
20'b00000101110000010110,
20'b00000110001011000001,
20'b00000101010110101100,
20'b00000101110000010110,
20'b00000101110100011101,
20'b00000101011101111000
};
#600;
reall[166] = 0;

pred [166] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 167 False
test_index = 16'd167;
x = {
20'b00000100101100011000,
20'b00000100110001010000,
20'b00000100110000000010,
20'b00000100110001010000,
20'b00000100100101000101,
20'b00000100100010101010,
20'b00000100100110010011,
20'b00000100011011010111,
20'b00000100011111000000,
20'b00000100101100011000
};
#600;
reall[167] = 0;

pred [167] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 168 False
test_index = 16'd168;
x = {
20'b00000011001101011010,
20'b00000100001001101101,
20'b00000100001101110010,
20'b00000100010100111100,
20'b00000100101101011110,
20'b00000011011010101100,
20'b00000011100101111100,
20'b00000100001100110001,
20'b00000011101110000111,
20'b00000011110011001110
};
#600;
reall[168] = 0;

pred [168] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 169 False
test_index = 16'd169;
x = {
20'b00000101010001100100,
20'b00000110010101010010,
20'b00000110001000111110,
20'b00000101100111000111,
20'b00000110000110111011,
20'b00000101111111101111,
20'b00000110010010001101,
20'b00000101101100001111,
20'b00000101011111111011,
20'b00000101111110101101
};
#600;
reall[169] = 0;

pred [169] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 170 True
test_index = 16'd170;
x = {
20'b00000101000000000000,
20'b00000100111101000001,
20'b00000100001000111011,
20'b00000011101011001010,
20'b00000110110001000111,
20'b00000011101001101011,
20'b00000110001011111010,
20'b00000101000001011111,
20'b00000011011001010011,
20'b00000110011101110001
};
#600;
reall[170] = 1;

pred [170] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 171 False
test_index = 16'd171;
x = {
20'b00000110011101011011,
20'b00000110011110110011,
20'b00000110100100010001,
20'b00000110010010011110,
20'b00000110011010101100,
20'b00000110011110110011,
20'b00000110011110110011,
20'b00000110010010011110,
20'b00000110010011110110,
20'b00000110010111111101
};
#600;
reall[171] = 0;

pred [171] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 172 False
test_index = 16'd172;
x = {
20'b00000101111101110010,
20'b00000101111000101110,
20'b00000101110100111100,
20'b00000101111101110010,
20'b00000101111000101110,
20'b00000101110001001001,
20'b00000101111000101110,
20'b00000101111011010000,
20'b00000110000110101000,
20'b00000110000010110110
};
#600;
reall[172] = 0;

pred [172] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 173 False
test_index = 16'd173;
x = {
20'b00000100110000001010,
20'b00000100110110011111,
20'b00000100101100010110,
20'b00000100101110111001,
20'b00000100101100010110,
20'b00000100110001011011,
20'b00000100101110111001,
20'b00000100110010101100,
20'b00000100110001011011,
20'b00000100101101100111
};
#600;
reall[173] = 0;

pred [173] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 174 False
test_index = 16'd174;
x = {
20'b00000101100010110000,
20'b00000101100111110010,
20'b00000101111101001010,
20'b00000110000000111100,
20'b00000101110100010111,
20'b00000101111101001010,
20'b00000101110100010111,
20'b00000101101001000010,
20'b00000101011110111110,
20'b00000101110011000110
};
#600;
reall[174] = 0;

pred [174] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 175 False
test_index = 16'd175;
x = {
20'b00000010000011100000,
20'b00000001100011100101,
20'b00000001101111000101,
20'b00000001101010110100,
20'b00000001100110100100,
20'b00000010000000111101,
20'b00000001001100100110,
20'b00000001001010011110,
20'b00000010110101010011,
20'b00000001110111100110
};
#600;
reall[175] = 0;

pred [175] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 176 False
test_index = 16'd176;
x = {
20'b00000110101001110000,
20'b00000110101101110111,
20'b00000110100000001010,
20'b00000110000111100001,
20'b00000101110101101110,
20'b00000101110111000110,
20'b00000101110100010111,
20'b00000110001110010111,
20'b00000110101100011111,
20'b00000110111100111010
};
#600;
reall[176] = 0;

pred [176] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 177 True
test_index = 16'd177;
x = {
20'b00000001110010001010,
20'b00000011011001000101,
20'b00000011011110010001,
20'b00000011001010011000,
20'b00000010111001111100,
20'b00000011100100010100,
20'b00000011000100010100,
20'b00000001110001010011,
20'b00000010111010110011,
20'b00000001111110010001
};
#600;
reall[177] = 1;

pred [177] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 178 True
test_index = 16'd178;
x = {
20'b00000101000000000000,
20'b00000011010000010111,
20'b00000110100000101111,
20'b00000101000100011101,
20'b00000101000100011101,
20'b00000011011001010011,
20'b00000110100101001101,
20'b00000101000010111110,
20'b00000100111000100011,
20'b00000011011001010011
};
#600;
reall[178] = 1;

pred [178] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 179 True
test_index = 16'd179;
x = {
20'b00000100101100101001,
20'b00000011010111110100,
20'b00000110000000000000,
20'b00000100110100000101,
20'b00000100111000100011,
20'b00000100101110001000,
20'b00000100101111101000,
20'b00000011010000010111,
20'b00000110000111011100,
20'b00000100101111101000
};
#600;
reall[179] = 1;

pred [179] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 180 True
test_index = 16'd180;
x = {
20'b00000100010110100101,
20'b00000011101001011010,
20'b00000010110100101101,
20'b00000101100101000110,
20'b00000011101111110111,
20'b00000011101000010101,
20'b00000011000101111010,
20'b00000100011101000010,
20'b00000011011000001100,
20'b00000100111001000000
};
#600;
reall[180] = 1;

pred [180] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 181 False
test_index = 16'd181;
x = {
20'b00000100110101000110,
20'b00000101000001110010,
20'b00000100110101000110,
20'b00000100111101000001,
20'b00000100111101000001,
20'b00000101000110100010,
20'b00000100110001111011,
20'b00000100111000010001,
20'b00000100111000010001,
20'b00000100111001110110
};
#600;
reall[181] = 0;

pred [181] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 182 False
test_index = 16'd182;
x = {
20'b00000100110110000111,
20'b00000100101110110100,
20'b00000100110011101011,
20'b00000100110111010101,
20'b00000101000011011111,
20'b00000101001001100100,
20'b00000101000111001001,
20'b00000100110110000111,
20'b00000100101001111101,
20'b00000100110100111001
};
#600;
reall[182] = 0;

pred [182] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 183 False
test_index = 16'd183;
x = {
20'b00000101000010010001,
20'b00000100111101011010,
20'b00000100110010011110,
20'b00000100100101000101,
20'b00000100101100011000,
20'b00000100110001010000,
20'b00000101000001000100,
20'b00000101000101111011,
20'b00000100111110101000,
20'b00000100111000100011
};
#600;
reall[183] = 0;

pred [183] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 184 False
test_index = 16'd184;
x = {
20'b00000110010001001100,
20'b00000110001101010111,
20'b00000110001001100011,
20'b00000110001001100011,
20'b00000110001111111010,
20'b00000110000001111010,
20'b00000101111010010001,
20'b00000110010010011101,
20'b00000110100000011110,
20'b00000110010010011101
};
#600;
reall[184] = 0;

pred [184] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 185 False
test_index = 16'd185;
x = {
20'b00000110000001111010,
20'b00000101110110011100,
20'b00000101101110110011,
20'b00000110001110101001,
20'b00000110011011011000,
20'b00000110010010011101,
20'b00000110010101000000,
20'b00000110001101010111,
20'b00000110001000010001,
20'b00000110000011001011
};
#600;
reall[185] = 0;

pred [185] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 186 False
test_index = 16'd186;
x = {
20'b00000101000000110010,
20'b00000101001101010111,
20'b00000101100100000000,
20'b00000101010011101001,
20'b00000101010001001000,
20'b00000101000000110010,
20'b00000101001001100101,
20'b00000101010010011001,
20'b00000101011011001101,
20'b00000101011000101100
};
#600;
reall[186] = 0;

pred [186] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 187 False
test_index = 16'd187;
x = {
20'b00000101110010010110,
20'b00000101111011001101,
20'b00000101101100011100,
20'b00000101101101111011,
20'b00000101111001101110,
20'b00000101101010111110,
20'b00000101111001101110,
20'b00000101101010111110,
20'b00000101110011110100,
20'b00000101101101111011
};
#600;
reall[187] = 0;

pred [187] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 188 False
test_index = 16'd188;
x = {
20'b00000110000111011011,
20'b00000110001100011000,
20'b00000110001110000010,
20'b00000110000100001000,
20'b00000110000100001000,
20'b00000110000100001000,
20'b00000101111000100100,
20'b00000101101110101010,
20'b00000101100110011001,
20'b00000110010010111111
};
#600;
reall[188] = 0;

pred [188] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 189 False
test_index = 16'd189;
x = {
20'b00000100100100101111,
20'b00000100011111111011,
20'b00000100011100010011,
20'b00000100100001001000,
20'b00000100101101001011,
20'b00000100100001001000,
20'b00000100011110101110,
20'b00000100011111111011,
20'b00000100100111001001,
20'b00000100100111001001
};
#600;
reall[189] = 0;

pred [189] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 190 False
test_index = 16'd190;
x = {
20'b00000111100101100001,
20'b00000111010011110111,
20'b00000111011100101100,
20'b00000111100110100111,
20'b00000111011101110010,
20'b00000111100100011010,
20'b00000111010010110000,
20'b00000111100110100111,
20'b00000111010010110000,
20'b00000111010111001011
};
#600;
reall[190] = 0;

pred [190] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 191 False
test_index = 16'd191;
x = {
20'b00000101100010011000,
20'b00000101010011001010,
20'b00000101011011110110,
20'b00000101010000111111,
20'b00000101010011001010,
20'b00000101010110011010,
20'b00000110000101001010,
20'b00000110000010111111,
20'b00000101010010000100,
20'b00000101111100011101
};
#600;
reall[191] = 0;

pred [191] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 192 False
test_index = 16'd192;
x = {
20'b00000101001100111000,
20'b00000100111110100111,
20'b00000100111000010001,
20'b00000101001000000111,
20'b00000101000011010111,
20'b00000101000000001100,
20'b00000101000000001100,
20'b00000101001001101101,
20'b00000101001001101101,
20'b00000100111101000001
};
#600;
reall[192] = 0;

pred [192] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 193 False
test_index = 16'd193;
x = {
20'b00000111001100001000,
20'b00000111010110000100,
20'b00000111011011100101,
20'b00000111010001101001,
20'b00000111100000000000,
20'b00000111001001111011,
20'b00000111010100111101,
20'b00000111000000000000,
20'b00000111010011110111,
20'b00000111010001101001
};
#600;
reall[193] = 0;

pred [193] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 194 False
test_index = 16'd194;
x = {
20'b00000100100000101101,
20'b00000100001000110100,
20'b00000100111101110010,
20'b00000100011110101000,
20'b00000100110001010101,
20'b00000100110110100001,
20'b00000100011100100011,
20'b00000100101011000110,
20'b00000100110001010101,
20'b00000100011101100110
};
#600;
reall[194] = 0;

pred [194] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 195 False
test_index = 16'd195;
x = {
20'b00000101011111000101,
20'b00000101100101111010,
20'b00000101101100101111,
20'b00000101100111110111,
20'b00000101101110101100,
20'b00000101101100101111,
20'b00000101101100101111,
20'b00000101110000101000,
20'b00000101101000110101,
20'b00000101101000110101
};
#600;
reall[195] = 0;

pred [195] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 196 False
test_index = 16'd196;
x = {
20'b00000100101000101110,
20'b00000101001110001000,
20'b00000101000011010100,
20'b00000100110110110110,
20'b00000100100111111001,
20'b00000100101011001110,
20'b00000100100111111001,
20'b00000101001000010011,
20'b00000110000110101001,
20'b00000100011101000101
};
#600;
reall[196] = 0;

pred [196] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 197 False
test_index = 16'd197;
x = {
20'b00000110011110110101,
20'b00000101110010111010,
20'b00000110000111011110,
20'b00000110001111111000,
20'b00000101110101101110,
20'b00000110001011001101,
20'b00000110001010010001,
20'b00000101110100110010,
20'b00000110110110001100,
20'b00000110001111111000
};
#600;
reall[197] = 0;

pred [197] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 198 True
test_index = 16'd198;
x = {
20'b00000000111111110010,
20'b00000000010011110100,
20'b00000001010011100111,
20'b00000100110111001010,
20'b00000010101101010000,
20'b00000100101001010111,
20'b00000010100011110001,
20'b00000010001000001100,
20'b00000000111101001100,
20'b00000011000101011000
};
#600;
reall[198] = 1;

pred [198] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 199 True
test_index = 16'd199;
x = {
20'b00000010000001110101,
20'b00000101011101000000,
20'b00000011111011011001,
20'b00000010001000010010,
20'b00000010111000001011,
20'b00000010111001000101,
20'b00000100001000010010,
20'b00000011110110110010,
20'b00000011100011011101,
20'b00000011100000101100
};
#600;
reall[199] = 1;

pred [199] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
        
        // Initialize variables
        sum = 0;
        true = 0;

        for (i = 0; i < max_data; i = i + 1) begin
            if (!(reall[i] === 1'bx || pred[i] === 1'bx)) begin
                $display("testcase: %d, real: %b, pred: %b", i, reall[i], pred[i]);
                sum = sum + 1;
                if (reall[i] == pred[i]) begin
                    true = true + 1;
                end
            end
        end

        if (sum > 0) begin
            $display("accuracy = (%d / %d) = %.3f%%", true, sum, true * 100.0 / sum);
        end else begin
            $display("No valid test cases to calculate accuracy.");
        end

        // Finish simulation
        $finish;
    end

    initial begin
        // // Initialize variables
        // sum = 0;
        // true = 0;

        // for (i = 0; i < 25; i = i + 1) begin
        //     if (!(reall[i] === 1'bx || pred[i] === 1'bx)) begin
        //         $display("testcase: %d, real: %b, pred: %b", i, reall[i], pred[i]);
        //         sum = sum + 1;
        //         if (reall[i] == pred[i]) begin
        //             true = true + 1;
        //         end
        //     end
        // end

        // if (sum > 0) begin
        //     $display("accuracy = %4d / %4d = %4f", true, sum, true * 1.0 / sum);
        // end else begin
        //     $display("No valid test cases to calculate accuracy.");
        // end
    end

endmodule
