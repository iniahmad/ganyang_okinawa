
`include "encoder_fixed_point.v"

`timescale 1ns / 1ps

module encoder_fixed_point_tb;
    // Parameters
    parameter N_input = 9;
    parameter M_output = 4;
    parameter BITSIZE = 32; // 1-bit sign, 4-bit exponent, 27-bit mantissa

    // Testbench signals
    reg [N_input * BITSIZE - 1:0] x;          // Input data
    reg [N_input * M_output * BITSIZE - 1:0] w; // Weights
    reg [M_output * BITSIZE - 1:0] b;         // Bias
    wire [M_output * BITSIZE - 1:0] out;      // Output data

    // Instantiate the DUT
    encoder_fixed_point #(
        .N_input(N_input),
        .M_output(M_output),
        .BITSIZE(BITSIZE)
    ) dut (
        .x(x),
        .w(w),
        .b(b),
        .out(out)
    );

    initial begin
        // $dumpfile("encoder_fixed_point_tb.vcd");
        // $dumpvars(0, encoder_fixed_point_tb);
        // Initialize inputs
        x = {
            32'b0_00101_0000000000000000000000001, // x[8] = 5.000001
            32'b0_00100_0000000000000000000000010, // x[7] = 4.000002
            32'b0_00011_0000000000000000000000011, // x[6] = 3.000003
            32'b0_00010_0000000000000000000000100, // x[5] = 2.000004
            32'b0_00001_0000000000000000000000101, // x[4] = 1.000005
            32'b0_00000_0000000000000000000000110, // x[3] = 0.000006
            32'b1_11111_0000000000000000000000111, // x[2] = -1.000007
            32'b1_11110_0000000000000000000001000, // x[1] = -2.000008
            32'b1_11101_0000000000000000000001001  // x[0] = -3.000009
        };

        w = {
            32'b0_00010_0000000000000000000001010, // w[35] = 2.00000A
            32'b0_00001_0000000000000000000001011, // w[34] = 1.00000B
            32'b0_00011_0000000000000000000001100, // ...
            32'b0_00000_0000000000000000000001101,
            32'b1_11111_0000000000000000000001110,
            32'b1_11110_0000000000000000000001111,
            32'b1_11101_0000000000000000000010000,
            32'b0_00100_0000000000000000000010001,
            32'b1_11100_0000000000000000000010010,
            32'b0_00101_0000000000000000000010011,
            32'b1_11101_0000000000000000000010100,
            32'b0_00000_0000000000000000000010101,
            32'b0_00001_0000000000000000000010110,
            32'b0_00010_0000000000000000000010111,
            32'b0_00011_0000000000000000000011000,
            32'b0_00100_0000000000000000000011001,
            32'b0_00010_0000000000000000000011010,
            32'b0_00001_0000000000000000000011011,
            32'b0_00011_0000000000000000000011100,
            32'b0_00000_0000000000000000000011101,
            32'b1_11111_0000000000000000000011110,
            32'b1_11110_0000000000000000000011111,
            32'b1_11101_0000000000000000000100000,
            32'b0_00100_0000000000000000000100001,
            32'b1_11100_0000000000000000000100010,
            32'b0_00101_0000000000000000000100011,
            32'b1_11101_0000000000000000000100100,
            32'b0_00000_0000000000000000000100101,
            32'b0_00001_0000000000000000000100110,
            32'b0_00010_0000000000000000000100111,
            32'b0_00011_0000000000000000000101000,
            32'b0_00100_0000000000000000000101001,
            32'b0_00011_0000000000000000000101010,
            32'b0_00001_0000000000000000000101011,
            32'b0_00010_0000000000000000000101100,
            32'b0_00000_0000000000000000000101101
        };

        b = {
            32'b0_00001_0000000000000000000100001, // b[3] = 1.000021
            32'b0_00010_0000000000000000000100010, // b[2] = 2.000022
            32'b0_00011_0000000000000000000100011, // b[1] = 3.000023
            32'b0_00100_0000000000000000000100100  // b[0] = 4.000024
        };

        // Wait for simulation
        #1000;

        // Display outputs
        $display("Output values:");
        $display("out[0] = %b", out[31:0]);
        $display("out[1] = %b", out[63:32]);
        $display("out[2] = %b", out[95:64]);
        $display("out[3] = %b", out[127:96]);

        // End simulation
        $stop;

    end
endmodule
