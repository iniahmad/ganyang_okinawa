`include "top_arrhythmia.v"

module top_arrhythmia_tb;

    // Parameters
    parameter BITSIZE = 24;

    // Inputs
    reg clk;
    reg reset;
    reg [BITSIZE*10-1:0] x;
    reg [6:0] test_index;
    // reg valid;

    // Outputs
    wire [BITSIZE-1:0] y1;
    wire [BITSIZE-1:0] y2;
    wire [BITSIZE*2-1:0] y;
    wire done_flag;
    // wire [BITSIZE-1:0] y2;

    // Instantiate the Unit Under Test (UUT)
    top_arrhythmia #(BITSIZE) uut (
        .clk(clk),
        .reset(reset),
        .x(x),
        .y({y1,y2}),
        .done_flag_out(done_flag)
    );

/// for output ///
    localparam max_data = 201;
    integer i;
    integer sum;
    integer true;
    logic pred  [max_data-1:0];
    logic reall [max_data-1:0];

    function logic compare_sign_mag;
        input [BITSIZE-1:0] val_a;
        input [BITSIZE-1:0] val_b;  // Declare inputs as 16-bit
        logic sign_a;
        logic sign_b;
        logic [BITSIZE-2:0] mag_a;
        logic [BITSIZE-2:0] mag_b;

        begin
            // Extract sign and magnitude
            sign_a = val_a[BITSIZE-1];
            sign_b = val_b[BITSIZE-1];
            mag_a = val_a[BITSIZE-2:0];
            mag_b = val_b[BITSIZE-2:0];

            // Compare based on sign and magnitude
            if (sign_a != sign_b) begin
                // If signs differ, the negative number is smaller
                compare_sign_mag = (sign_a < sign_b);  // 1 if A > B
            end else begin
                // If signs are the same, compare magnitudes
                if (sign_a == 1'b1) begin
                    // Both negative: larger magnitude means smaller number
                    compare_sign_mag = (mag_a < mag_b);  // 1 if (-)A > (-)B
                end else begin
                    // Both positive: larger magnitude means larger number
                    compare_sign_mag = (mag_a > mag_b);  // 1 if A > B
                end
            end
        end
    endfunction
/// for output ///

    // Clock generation
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 10 time units period
    end

    // Test sequence
    initial begin
        // $dumpfile("top_arrhythmia_tb.vcd");
        // $dumpvars(0, top_arrhythmia_tb);
        // Initialize Inputs
        reset = 1;
        x = 0;

        // Wait for global reset to finish
        #10;
        reset = 0;

// Testcase 0 True
test_index = 16'd0;
x = {
24'b000000000100001011000011,
24'b000000000001111111000101,
24'b000000000110010111111100,
24'b000000000100011001110010,
24'b000000000100001101110100,
24'b000000000001010011110011,
24'b000000000001010100101110,
24'b000000000101111010011110,
24'b000000000011101101100101,
24'b000000000010101111111000
};
#600;
reall[0] = 1;

pred [0] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 1 False
test_index = 16'd1;
x = {
24'b000000000100011100011100,
24'b000000000011101101000010,
24'b000000000011010010010100,
24'b000000000011011010111011,
24'b000000000010101011100001,
24'b000000000100100110110010,
24'b000000000010101001110011,
24'b000000000100001100000100,
24'b000000000011100110001001,
24'b000000000011011010111011
};
#600;
reall[1] = 0;

pred [1] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 2 False
test_index = 16'd2;
x = {
24'b000000000101110110111000,
24'b000000000110000011011101,
24'b000000000101111110011011,
24'b000000000101110100010111,
24'b000000000101101011100011,
24'b000000000101101010010011,
24'b000000000101100001011111,
24'b000000000101101110000100,
24'b000000000101110011000110,
24'b000000000110000010001100
};
#600;
reall[2] = 0;

pred [2] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 3 True
test_index = 16'd3;
x = {
24'b000000000011010101000100,
24'b000000000010110110010001,
24'b000000000010111010010101,
24'b000000000011001011010101,
24'b000000000010110100101010,
24'b000000000010111001100001,
24'b000000000011000011001111,
24'b000000000010001100111101,
24'b000000000100010111011111,
24'b000000000011010001110100
};
#600;
reall[3] = 1;

pred [3] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 4 True
test_index = 16'd4;
x = {
24'b000000000011101110110010,
24'b000000000110010111101010,
24'b000000000010111010000101,
24'b000000000101101111110111,
24'b000000000011010110000011,
24'b000000000011000010101100,
24'b000000000011000010101100,
24'b000000000100101110010000,
24'b000000000100100101101001,
24'b000000000100110101110010
};
#600;
reall[4] = 1;

pred [4] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 5 False
test_index = 16'd5;
x = {
24'b000000000101100110100001,
24'b000000000101010010011001,
24'b000000000101010110001011,
24'b000000000101111101001010,
24'b000000000110000000111100,
24'b000000000101011110111110,
24'b000000000101100100000000,
24'b000000000101100110100001,
24'b000000000101101011100011,
24'b000000000101010001001000
};
#600;
reall[5] = 0;

pred [5] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 6 True
test_index = 16'd6;
x = {
24'b000000000100011000111100,
24'b000000000010101111111010,
24'b000000001000000000000000,
24'b000000000101111011011001,
24'b000000000101110011100001,
24'b000000000011110000001111,
24'b000000000111100101101111,
24'b000000000101111011011001,
24'b000000000101110111011101,
24'b000000000011101101100111
};
#600;
reall[6] = 1;

pred [6] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 7 True
test_index = 16'd7;
x = {
24'b000000000100010110100101,
24'b000000000011110110010100,
24'b000000000011001011010010,
24'b000000000100100110101110,
24'b000000000001110010000001,
24'b000000000001110011000101,
24'b000000000111010010110100,
24'b000000000011010110000011,
24'b000000000101101101101101,
24'b000000000011100010111101
};
#600;
reall[7] = 1;

pred [7] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 8 False
test_index = 16'd8;
x = {
24'b000000000110010001000111,
24'b000000000110010001000111,
24'b000000000101100001010010,
24'b000000000101011111000111,
24'b000000000101111100011101,
24'b000000000110000000110100,
24'b000000000101111000000111,
24'b000000000101010110011010,
24'b000000000101111110101001,
24'b000000000110010011010010
};
#600;
reall[8] = 0;

pred [8] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 9 False
test_index = 16'd9;
x = {
24'b000000000110000011111110,
24'b000000000101111010011011,
24'b000000000101110000111001,
24'b000000000110001011111011,
24'b000000000110000111001001,
24'b000000000101111111001101,
24'b000000000101110101101010,
24'b000000000101111111001101,
24'b000000000101111000110110,
24'b000000000110000011111110
};
#600;
reall[9] = 0;

pred [9] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 10 True
test_index = 16'd10;
x = {
24'b000000000001011111011100,
24'b000000000010000110110111,
24'b000000000001110110010001,
24'b000000000001110001000101,
24'b000000000001101000010001,
24'b000000000010101000000100,
24'b000000000001100111101111,
24'b000000000010000110110111,
24'b000000000001110100001100,
24'b000000000001100101001001
};
#600;
reall[10] = 1;

pred [10] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 11 True
test_index = 16'd11;
x = {
24'b000000000010111101100100,
24'b000000000011000100110111,
24'b000000000001000110011110,
24'b000000000001000110011110,
24'b000000000100010010101000,
24'b000000000011010111011111,
24'b000000000001010011011100,
24'b000000000000110011110110,
24'b000000000011100010110101,
24'b000000000011110010001110
};
#600;
reall[11] = 1;

pred [11] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 12 False
test_index = 16'd12;
x = {
24'b000000000101111111101000,
24'b000000000101111110001001,
24'b000000000101111011001101,
24'b000000000101111100101011,
24'b000000000110001011011011,
24'b000000000101111011001101,
24'b000000000110000001000110,
24'b000000000101110110110001,
24'b000000000101110101010011,
24'b000000000101111011001101
};
#600;
reall[12] = 0;

pred [12] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 13 False
test_index = 16'd13;
x = {
24'b000000000100111011101101,
24'b000000000101000000111010,
24'b000000000100111100110000,
24'b000000000101000000111010,
24'b000000000100111110110101,
24'b000000000100111111110111,
24'b000000000101001100010101,
24'b000000000100011100100011,
24'b000000000101011011111010,
24'b000000000101001111011100
};
#600;
reall[13] = 0;

pred [13] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 14 True
test_index = 16'd14;
x = {
24'b000000000011000000110111,
24'b000000000101100000000000,
24'b000000000010111100100010,
24'b000000000101000110111010,
24'b000000000011110011111001,
24'b000000000011100000110111,
24'b000000000011110101100111,
24'b000000000100101101110101,
24'b000000000100011001000101,
24'b000000000100011100100010
};
#600;
reall[14] = 1;

pred [14] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 15 False
test_index = 16'd15;
x = {
24'b000000000101101111010011,
24'b000000000101101000111100,
24'b000000000101101100000111,
24'b000000000101100010100101,
24'b000000000101110000111001,
24'b000000000101110010011111,
24'b000000000101101100000111,
24'b000000000101100010100101,
24'b000000000101101000111100,
24'b000000000101101010100010
};
#600;
reall[15] = 0;

pred [15] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 16 True
test_index = 16'd16;
x = {
24'b000000000110001101011001,
24'b000000000100111010000010,
24'b000000000100101111101000,
24'b000000000100110100000101,
24'b000000000100101110001000,
24'b000000000100110001000111,
24'b000000000011000111011100,
24'b000000000110011001010011,
24'b000000000100011010110010,
24'b000000000101001010011010
};
#600;
reall[16] = 1;

pred [16] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 17 False
test_index = 16'd17;
x = {
24'b000000000101110011011010,
24'b000000000101111010010110,
24'b000000000101101101010101,
24'b000000000101011011000111,
24'b000000000101011101101110,
24'b000000000101101111111100,
24'b000000000101110111110000,
24'b000000000101100110011001,
24'b000000000101010111101001,
24'b000000000101011100110110
};
#600;
reall[17] = 0;

pred [17] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 18 False
test_index = 16'd18;
x = {
24'b000000000010110010001110,
24'b000000000011001100111101,
24'b000000000010111111001100,
24'b000000000010110110010001,
24'b000000000010111100110000,
24'b000000000011101011101111,
24'b000000000011010111011111,
24'b000000000100001101110001,
24'b000000000010101110001011,
24'b000000000010110100101010
};
#600;
reall[18] = 0;

pred [18] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 19 False
test_index = 16'd19;
x = {
24'b000000000101100100000000,
24'b000000000101100101010001,
24'b000000000101110100010111,
24'b000000000101111001011001,
24'b000000000101111110011011,
24'b000000000101101100110100,
24'b000000000101100001011111,
24'b000000000101100000001111,
24'b000000000101100100000000,
24'b000000000101101110000100
};
#600;
reall[19] = 0;

pred [19] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 20 False
test_index = 16'd20;
x = {
24'b000000000100111000100001,
24'b000000000100101111011000,
24'b000000000100111011110110,
24'b000000000100111100101011,
24'b000000000100101011001110,
24'b000000000100111011000000,
24'b000000000100110100010111,
24'b000000000111001101010011,
24'b000000000011101100111000,
24'b000000000101011011011011
};
#600;
reall[20] = 0;

pred [20] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 21 False
test_index = 16'd21;
x = {
24'b000000000101100000001110,
24'b000000000101011110010111,
24'b000000000110011011000110,
24'b000000000110110100010100,
24'b000000000110100111001111,
24'b000000000111001001110011,
24'b000000000110110100010100,
24'b000000000101110011110110,
24'b000000000110010111010110,
24'b000000000110010110011011
};
#600;
reall[21] = 0;

pred [21] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 22 False
test_index = 16'd22;
x = {
24'b000000000011010100111001,
24'b000000000011010010010100,
24'b000000000100011011100101,
24'b000000000011101010011100,
24'b000000000011100101010001,
24'b000000000100000100010011,
24'b000000000100110000010001,
24'b000000000101000100000110,
24'b000000000011100011100011,
24'b000000000011100101010001
};
#600;
reall[22] = 0;

pred [22] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 23 False
test_index = 16'd23;
x = {
24'b000000000101111111001011,
24'b000000000101111010001110,
24'b000000000101011001001011,
24'b000000000110010111111100,
24'b000000000101101110101010,
24'b000000000110001010101111,
24'b000000000110011001100110,
24'b000000000110010100101001,
24'b000000000110000100001000,
24'b000000000101111111001011
};
#600;
reall[23] = 0;

pred [23] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 24 False
test_index = 16'd24;
x = {
24'b000000000110000101100010,
24'b000000000110000010100101,
24'b000000000110000010100101,
24'b000000000110001110011000,
24'b000000000110001001111101,
24'b000000000110000101100010,
24'b000000000110001000011110,
24'b000000000110010100010010,
24'b000000000110010001010101,
24'b000000000101111110001001
};
#600;
reall[24] = 0;

pred [24] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 25 False
test_index = 16'd25;
x = {
24'b000000000100100111000011,
24'b000000000100011110010111,
24'b000000000100000111001110,
24'b000000000100001000101011,
24'b000000000100001011100100,
24'b000000000100000100010101,
24'b000000000100001101000001,
24'b000000000100001101000001,
24'b000000000100100001010000,
24'b000000000011101011110000
};
#600;
reall[25] = 0;

pred [25] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 26 False
test_index = 16'd26;
x = {
24'b000000000100011011011110,
24'b000000000100011111110100,
24'b000000000100100100001010,
24'b000000000100101011011000,
24'b000000000100100100001010,
24'b000000000100011011011110,
24'b000000000100001111111010,
24'b000000000100001010000111,
24'b000000000100001011100100,
24'b000000000100010100001111
};
#600;
reall[26] = 0;

pred [26] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 27 False
test_index = 16'd27;
x = {
24'b000000000010101010001000,
24'b000000000011110001011010,
24'b000000000011000100110111,
24'b000000000011111000101101,
24'b000000000010101100100011,
24'b000000000010101010001000,
24'b000000000010100001001101,
24'b000000000010101011101111,
24'b000000000011001000111010,
24'b000000000011011101111110
};
#600;
reall[27] = 0;

pred [27] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 28 True
test_index = 16'd28;
x = {
24'b000000000101000010111110,
24'b000000000100110101100101,
24'b000000000100111000100011,
24'b000000000100101100101001,
24'b000000000100111000100011,
24'b000000000100011010110010,
24'b000000000101010011010110,
24'b000000000100111110100000,
24'b000000000011010100110101,
24'b000000000110011001010011
};
#600;
reall[28] = 1;

pred [28] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 29 False
test_index = 16'd29;
x = {
24'b000000000101111000110110,
24'b000000000110000000110010,
24'b000000000110000111001001,
24'b000000000101111010011011,
24'b000000000101110101101010,
24'b000000000101111101100111,
24'b000000000110001000101111,
24'b000000000101111010011011,
24'b000000000101101100000111,
24'b000000000101110000111001
};
#600;
reall[29] = 0;

pred [29] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 30 True
test_index = 16'd30;
x = {
24'b000000000110000110110111,
24'b000000000010111000100011,
24'b000000000010101011010011,
24'b000000000011011001101010,
24'b000000000011000101110010,
24'b000000000100011010111110,
24'b000000000100100011011111,
24'b000000000101001000011001,
24'b000000000011000100110110,
24'b000000000111001100111001
};
#600;
reall[30] = 1;

pred [30] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 31 True
test_index = 16'd31;
x = {
24'b000000000001100101001100,
24'b000000000011001100000110,
24'b000000000001110100110000,
24'b000000000100010010001010,
24'b000000000011111110010001,
24'b000000000010001011001111,
24'b000000000011011000001101,
24'b000000000011110011111001,
24'b000000000010100000000000,
24'b000000000011001000101001
};
#600;
reall[31] = 1;

pred [31] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 32 False
test_index = 16'd32;
x = {
24'b000000000100110101110111,
24'b000000000101001110011111,
24'b000000000101100000111101,
24'b000000000101101100001111,
24'b000000000101010110101100,
24'b000000000101010110101100,
24'b000000000101010111101110,
24'b000000000101000111010011,
24'b000000000100110001110000,
24'b000000000101000101010000
};
#600;
reall[32] = 0;

pred [32] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 33 False
test_index = 16'd33;
x = {
24'b000000000110100100001011,
24'b000000000110100001000100,
24'b000000000110100100001011,
24'b000000000110101000110110,
24'b000000000110110110110110,
24'b000000000111000000001100,
24'b000000000110111101000101,
24'b000000000110110010001100,
24'b000000000110111110101000,
24'b000000000111000111111110
};
#600;
reall[33] = 0;

pred [33] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 34 False
test_index = 16'd34;
x = {
24'b000000000101011001110001,
24'b000000000101100111000111,
24'b000000000110001101000101,
24'b000000000101011110111010,
24'b000000000101011110111010,
24'b000000000101111101101100,
24'b000000000110111011010000,
24'b000000000101111000100011,
24'b000000000101110010011001,
24'b000000000110001011000001
};
#600;
reall[34] = 0;

pred [34] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 35 False
test_index = 16'd35;
x = {
24'b000000000101110010011111,
24'b000000000101111111001101,
24'b000000000110000101100100,
24'b000000000101111100000001,
24'b000000000101110010011111,
24'b000000000101110111010000,
24'b000000000101111000110110,
24'b000000000110000011111110,
24'b000000000110001000101111,
24'b000000000101110101101010
};
#600;
reall[35] = 0;

pred [35] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 36 True
test_index = 16'd36;
x = {
24'b000000000100111010011011,
24'b000000000001011101111101,
24'b000000000010100001011011,
24'b000000000101100111000000,
24'b000000000100010000010000,
24'b000000000101011101010111,
24'b000000000100011111111011,
24'b000000000100111100110101,
24'b000000000100011100010011,
24'b000000000101000000011100
};
#600;
reall[36] = 1;

pred [36] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 37 False
test_index = 16'd37;
x = {
24'b000000000100111000011010,
24'b000000000100011111110100,
24'b000000000100011000100101,
24'b000000000100000111001110,
24'b000000000100000101110010,
24'b000000000100001000101011,
24'b000000000100010010110011,
24'b000000000100011100111011,
24'b000000000100100111000011,
24'b000000000100110100000100
};
#600;
reall[37] = 0;

pred [37] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 38 True
test_index = 16'd38;
x = {
24'b000000000010101100001111,
24'b000000000010101111000101,
24'b000000000110000100111101,
24'b000000000010010101100001,
24'b000000000101110100111000,
24'b000000000010100110100100,
24'b000000000101110011111011,
24'b000000000010111111001011,
24'b000000000101100010111001,
24'b000000000010110001111011
};
#600;
reall[38] = 1;

pred [38] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 39 False
test_index = 16'd39;
x = {
24'b000000000100110010101100,
24'b000000000100110011111101,
24'b000000000100101110111001,
24'b000000000100101001110100,
24'b000000000100101110111001,
24'b000000000100111001000001,
24'b000000000100101100010110,
24'b000000000100101011000101,
24'b000000000100101001110100,
24'b000000000100110001011011
};
#600;
reall[39] = 0;

pred [39] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 40 False
test_index = 16'd40;
x = {
24'b000000000110001111111100,
24'b000000000110001001101110,
24'b000000000110000001111100,
24'b000000000110010100100111,
24'b000000000110010011000100,
24'b000000000110001111111100,
24'b000000000110000110100111,
24'b000000000110010011000100,
24'b000000000110001110011001,
24'b000000000110001111111100
};
#600;
reall[40] = 0;

pred [40] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 41 False
test_index = 16'd41;
x = {
24'b000000000101101100001111,
24'b000000000101111011101000,
24'b000000000110000000110001,
24'b000000000101111011101000,
24'b000000000101011010110011,
24'b000000000110010000001010,
24'b000000000110100110101110,
24'b000000000110000111111100,
24'b000000000101000010001011,
24'b000000000101000011001101
};
#600;
reall[41] = 0;

pred [41] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 42 False
test_index = 16'd42;
x = {
24'b000000000101101101010001,
24'b000000000110000011110110,
24'b000000000110000111111100,
24'b000000000101011100110110,
24'b000000000100111000111100,
24'b000000000101100101000100,
24'b000000000110010010001101,
24'b000000000110011101011111,
24'b000000000101110100011101,
24'b000000000101111100101010
};
#600;
reall[42] = 0;

pred [42] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 43 True
test_index = 16'd43;
x = {
24'b000000000010111011011010,
24'b000000000111001110101110,
24'b000000000010111100011000,
24'b000000000111001001111001,
24'b000000000010111010011100,
24'b000000000111010000101010,
24'b000000000010111100011000,
24'b000000000011100010000011,
24'b000000000011100011000001,
24'b000000000100111011111001
};
#600;
reall[43] = 1;

pred [43] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 44 False
test_index = 16'd44;
x = {
24'b000000000101100011110001,
24'b000000000101101011101001,
24'b000000000101101100111101,
24'b000000000101100110011001,
24'b000000000101101001000001,
24'b000000000101101110010001,
24'b000000000101100011110001,
24'b000000000101101001000001,
24'b000000000101011110100001,
24'b000000000101011101001101
};
#600;
reall[44] = 0;

pred [44] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 45 False
test_index = 16'd45;
x = {
24'b000000000111010000100011,
24'b000000000111001000110100,
24'b000000000111011001011000,
24'b000000000111010111001011,
24'b000000000111001011000010,
24'b000000000111011101110010,
24'b000000000111001011000010,
24'b000000000111010010110000,
24'b000000000111000111101110,
24'b000000000111010000100011
};
#600;
reall[45] = 0;

pred [45] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 46 False
test_index = 16'd46;
x = {
24'b000000000110000001111010,
24'b000000000110000101101110,
24'b000000000110010111100011,
24'b000000000110101010101010,
24'b000000000110101001011001,
24'b000000000110010001001100,
24'b000000000110000111000000,
24'b000000000110010110010010,
24'b000000000110100110110110,
24'b000000000110100110110110
};
#600;
reall[46] = 0;

pred [46] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 47 True
test_index = 16'd47;
x = {
24'b000000000111110101100101,
24'b000000000110010011001010,
24'b000000000010110010110111,
24'b000000000010100001110101,
24'b000000000111011010001001,
24'b000000000110011001110010,
24'b000000000011000001000100,
24'b000000000010101101001100,
24'b000000000111101001010010,
24'b000000000110001001101100
};
#600;
reall[47] = 1;

pred [47] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 48 False
test_index = 16'd48;
x = {
24'b000000000100110101001001,
24'b000000000100111010000001,
24'b000000000100110011001100,
24'b000000000100101100010111,
24'b000000000100110001001111,
24'b000000000100110111000110,
24'b000000000100101001011100,
24'b000000000100100110100001,
24'b000000000100101111010011,
24'b000000000100101001011100
};
#600;
reall[48] = 0;

pred [48] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 49 False
test_index = 16'd49;
x = {
24'b000000000011010101011110,
24'b000000000011000100000111,
24'b000000000010100000100010,
24'b000000000011110101100101,
24'b000000000011111001111011,
24'b000000000100000110000100,
24'b000000000010011001100110,
24'b000000000100000110111100,
24'b000000000010001111001011,
24'b000000000100010100110100
};
#600;
reall[49] = 0;

pred [49] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 50 True
test_index = 16'd50;
x = {
24'b000000000111000110111111,
24'b000000000011111000011110,
24'b000000000101110010000001,
24'b000000000011101011100100,
24'b000000000100100011011111,
24'b000000000011000001100111,
24'b000000000101011000001100,
24'b000000000011101000010101,
24'b000000000100111011001010,
24'b000000000011100111010000
};
#600;
reall[50] = 1;

pred [50] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 51 True
test_index = 16'd51;
x = {
24'b000000000001101111100100,
24'b000000000011010101100111,
24'b000000000011011011101011,
24'b000000000011011001000101,
24'b000000000010000000110111,
24'b000000000101110011000001,
24'b000000000010000001101110,
24'b000000000011101101110101,
24'b000000000011011001111100,
24'b000000000011000000000000
};
#600;
reall[51] = 1;

pred [51] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 52 False
test_index = 16'd52;
x = {
24'b000000000110010111100011,
24'b000000000110000101101110,
24'b000000000110001100000110,
24'b000000000110001000010001,
24'b000000000110100001110000,
24'b000000000110011101111011,
24'b000000000110101010101010,
24'b000000000110100101100100,
24'b000000000110000101101110,
24'b000000000110001101010111
};
#600;
reall[52] = 0;

pred [52] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 53 True
test_index = 16'd53;
x = {
24'b000000000011110000111100,
24'b000000000100001100111010,
24'b000000000001101000010101,
24'b000000000001101000010101,
24'b000000000100011001110100,
24'b000000000011001101011100,
24'b000000000100110010100011,
24'b000000000011001101011100,
24'b000000000100110010100011,
24'b000000000011011101100101
};
#600;
reall[53] = 1;

pred [53] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 54 False
test_index = 16'd54;
x = {
24'b000000000010100011001001,
24'b000000000011110101100101,
24'b000000000011011111000001,
24'b000000000101000111001010,
24'b000000000010110000001010,
24'b000000000010110000001010,
24'b000000000010101010111101,
24'b000000000010111011011100,
24'b000000000011101110101001,
24'b000000000010111110111010
};
#600;
reall[54] = 0;

pred [54] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 55 False
test_index = 16'd55;
x = {
24'b000000000100100100101111,
24'b000000000100111011101000,
24'b000000000100100100101111,
24'b000000000100100100101111,
24'b000000000100100001001000,
24'b000000000100101001100011,
24'b000000000100100101111100,
24'b000000000100101001100011,
24'b000000000100100100101111,
24'b000000000100100100101111
};
#600;
reall[55] = 0;

pred [55] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 56 False
test_index = 16'd56;
x = {
24'b000000000101110101101010,
24'b000000000101101111010011,
24'b000000000101101100000111,
24'b000000000101100100001011,
24'b000000000101101010100010,
24'b000000000101100111010110,
24'b000000000101110010011111,
24'b000000000101111000110110,
24'b000000000101100111010110,
24'b000000000101100100001011
};
#600;
reall[56] = 0;

pred [56] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 57 False
test_index = 16'd57;
x = {
24'b000000000100100110000001,
24'b000000000100101011000101,
24'b000000000100100111010010,
24'b000000000100110001011011,
24'b000000000100110010101100,
24'b000000000100101101100111,
24'b000000000100100010001101,
24'b000000000100100111010010,
24'b000000000100101101100111,
24'b000000000100101101100111
};
#600;
reall[57] = 0;

pred [57] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 58 False
test_index = 16'd58;
x = {
24'b000000000101110111010000,
24'b000000000101111010011011,
24'b000000000110000000110010,
24'b000000000110000011111110,
24'b000000000110000011111110,
24'b000000000101111100000001,
24'b000000000101111000110110,
24'b000000000101111101100111,
24'b000000000110001011111011,
24'b000000000110000000110010
};
#600;
reall[58] = 0;

pred [58] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 59 False
test_index = 16'd59;
x = {
24'b000000000101110010101011,
24'b000000000110101001000010,
24'b000000000101101110010101,
24'b000000000101100011011101,
24'b000000000110001100110001,
24'b000000000110000010111111,
24'b000000000101011001101011,
24'b000000000101000011111100,
24'b000000000101110001100110,
24'b000000000101101101001111
};
#600;
reall[59] = 0;

pred [59] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 60 True
test_index = 16'd60;
x = {
24'b000000000001110101100111,
24'b000000000001101100111110,
24'b000000000011101001100000,
24'b000000000010000101001100,
24'b000000000010100111110010,
24'b000000000010111101011001,
24'b000000000010111011101011,
24'b000000000011010110011111,
24'b000000000010001111100100,
24'b000000000010001000101001
};
#600;
reall[60] = 1;

pred [60] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 61 True
test_index = 16'd61;
x = {
24'b000000000100000111101001,
24'b000000000010000100101011,
24'b000000000100010101010000,
24'b000000000010000001010001,
24'b000000000100010000001010,
24'b000000000001111011000010,
24'b000000000100010000001010,
24'b000000000010000110111100,
24'b000000000100010101110101,
24'b000000000001111111000000
};
#600;
reall[61] = 1;

pred [61] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 62 False
test_index = 16'd62;
x = {
24'b000000000101001111111001,
24'b000000000101011000100110,
24'b000000000101100010011000,
24'b000000000101011010110001,
24'b000000000101110010101011,
24'b000000000111000110011000,
24'b000000000110011011111111,
24'b000000000110010101011110,
24'b000000000110000010111111,
24'b000000000101110001100110
};
#600;
reall[62] = 0;

pred [62] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 63 False
test_index = 16'd63;
x = {
24'b000000000011001110110111,
24'b000000000011110011000100,
24'b000000000100010000011000,
24'b000000000100010000011000,
24'b000000000100001110101001,
24'b000000000100011100011100,
24'b000000000011010110101000,
24'b000000000011101101000010,
24'b000000000011001000110101,
24'b000000000011111111001000
};
#600;
reall[63] = 0;

pred [63] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 64 False
test_index = 16'd64;
x = {
24'b000000000101101010010011,
24'b000000000101101001000010,
24'b000000000101100000001111,
24'b000000000101111110011011,
24'b000000000110000111001110,
24'b000000000101011101101110,
24'b000000000101010100111010,
24'b000000000101100110100001,
24'b000000000101110001110110,
24'b000000000101110000100101
};
#600;
reall[64] = 0;

pred [64] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 65 False
test_index = 16'd65;
x = {
24'b000000000101110000010011,
24'b000000000101110000010011,
24'b000000000101100100101111,
24'b000000000101110110111010,
24'b000000000110001110000010,
24'b000000000110010010111111,
24'b000000000110000000110100,
24'b000000000101110110111010,
24'b000000000101111000100100,
24'b000000000101111011110111
};
#600;
reall[65] = 0;

pred [65] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 66 False
test_index = 16'd66;
x = {
24'b000000000110000001000110,
24'b000000000101111000010000,
24'b000000000110001001111101,
24'b000000000101111100101011,
24'b000000000110000101100010,
24'b000000000110001100111010,
24'b000000000110000101100010,
24'b000000000110000101100010,
24'b000000000110001111110111,
24'b000000000110001011011011
};
#600;
reall[66] = 0;

pred [66] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 67 False
test_index = 16'd67;
x = {
24'b000000000100100100011011,
24'b000000000100111110111011,
24'b000000000101000110100000,
24'b000000000100110011100101,
24'b000000000100100011011111,
24'b000000000100100111010001,
24'b000000000100101110110110,
24'b000000000101000000110100,
24'b000000000101010100101100,
24'b000000000101010100101100
};
#600;
reall[67] = 0;

pred [67] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 68 False
test_index = 16'd68;
x = {
24'b000000000110010100010000,
24'b000000000101110011011011,
24'b000000000101010001100100,
24'b000000000110010101010010,
24'b000000000110001000111110,
24'b000000000101100111000111,
24'b000000000110000110111011,
24'b000000000101111111101111,
24'b000000000110010010001101,
24'b000000000101101100001111
};
#600;
reall[68] = 0;

pred [68] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 69 False
test_index = 16'd69;
x = {
24'b000000000110001010111000,
24'b000000000110000101010011,
24'b000000000110011110111101,
24'b000000000110100011011010,
24'b000000000110011001011000,
24'b000000000110010010101011,
24'b000000000110001010111000,
24'b000000000110001000101001,
24'b000000000110010011110011,
24'b000000000110110100001001
};
#600;
reall[69] = 0;

pred [69] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 70 True
test_index = 16'd70;
x = {
24'b000000000001111001011000,
24'b000000000001110100101101,
24'b000000000001011110011010,
24'b000000000010000110110111,
24'b000000000001100111101111,
24'b000000000001101100011010,
24'b000000000001101111100001,
24'b000000000001101101111110,
24'b000000000010000100110011,
24'b000000000001110011101011
};
#600;
reall[70] = 1;

pred [70] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 71 False
test_index = 16'd71;
x = {
24'b000000000100001010111001,
24'b000000000010100100000101,
24'b000000000010011101110110,
24'b000000000010110000100011,
24'b000000000010101011010110,
24'b000000000010010111101000,
24'b000000000011101000101000,
24'b000000000010111000110111,
24'b000000000011000001001010,
24'b000000000011011111010010
};
#600;
reall[71] = 0;

pred [71] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 72 False
test_index = 16'd72;
x = {
24'b000000000100001011100100,
24'b000000000100100001010000,
24'b000000000100011000100101,
24'b000000000100101011011000,
24'b000000000100100101100110,
24'b000000000100100101100110,
24'b000000000100000111001110,
24'b000000000100001011100100,
24'b000000000100000010111001,
24'b000000000100001101000001
};
#600;
reall[72] = 0;

pred [72] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 73 False
test_index = 16'd73;
x = {
24'b000000000110011101011011,
24'b000000000110100001100010,
24'b000000000110111010001011,
24'b000000000110111010001011,
24'b000000000110111000110100,
24'b000000000110010101001110,
24'b000000000110000110001010,
24'b000000000101111101111100,
24'b000000000110001101000000,
24'b000000000110101101110111
};
#600;
reall[73] = 0;

pred [73] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 74 False
test_index = 16'd74;
x = {
24'b000000000101101100000111,
24'b000000000101110100000100,
24'b000000000101101111010011,
24'b000000000101111100000001,
24'b000000000101110111010000,
24'b000000000101110111010000,
24'b000000000101101010100010,
24'b000000000101111111001101,
24'b000000000101111010011011,
24'b000000000101110101101010
};
#600;
reall[74] = 0;

pred [74] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 75 False
test_index = 16'd75;
x = {
24'b000000000110110000110011,
24'b000000000110110101010000,
24'b000000000110010011110011,
24'b000000000110011011100110,
24'b000000000110010100111010,
24'b000000000110010110000001,
24'b000000000110100010010011,
24'b000000000110110100001001,
24'b000000000110101010000110,
24'b000000000110001011111111
};
#600;
reall[75] = 0;

pred [75] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 76 False
test_index = 16'd76;
x = {
24'b000000000110010011000100,
24'b000000000110100001000100,
24'b000000000110010111101110,
24'b000000000110011010110110,
24'b000000000110011111100000,
24'b000000000110101010011010,
24'b000000000110011001010010,
24'b000000000110011100011001,
24'b000000000110011111100000,
24'b000000000110011111100000
};
#600;
reall[76] = 0;

pred [76] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 77 False
test_index = 16'd77;
x = {
24'b000000000100110101001000,
24'b000000000100110011001100,
24'b000000000100110110000110,
24'b000000000100111000111111,
24'b000000000100110001010001,
24'b000000000100101101011001,
24'b000000000100111001111101,
24'b000000000100111000111111,
24'b000000000100110000010011,
24'b000000000100111001111101
};
#600;
reall[77] = 0;

pred [77] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 78 False
test_index = 16'd78;
x = {
24'b000000000100100111001001,
24'b000000000100101000010110,
24'b000000000100110001111111,
24'b000000000100101010110001,
24'b000000000100100011100010,
24'b000000000100011110101110,
24'b000000000100101001100011,
24'b000000000100101001100011,
24'b000000000100101010110001,
24'b000000000011010000011010
};
#600;
reall[78] = 0;

pred [78] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 79 True
test_index = 16'd79;
x = {
24'b000000000001101001010011,
24'b000000000010000111011001,
24'b000000000001110100001100,
24'b000000000001101010010101,
24'b000000000001001010001011,
24'b000000000001001010001011,
24'b000000000001110101001111,
24'b000000000001011110011010,
24'b000000000001011011110100,
24'b000000000010011101101100
};
#600;
reall[79] = 1;

pred [79] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 80 False
test_index = 16'd80;
x = {
24'b000000000101001111111001,
24'b000000000101101000111001,
24'b000000000101111101100011,
24'b000000000101001111111001,
24'b000000000100111110100000,
24'b000000000101001100101000,
24'b000000000101001110110011,
24'b000000000101001100101000,
24'b000000000100111100010101,
24'b000000000101000010110110
};
#600;
reall[80] = 0;

pred [80] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 81 False
test_index = 16'd81;
x = {
24'b000000000101100100000000,
24'b000000000101100110100001,
24'b000000000101101011100011,
24'b000000000101010001001000,
24'b000000000101011100011101,
24'b000000000101101010010011,
24'b000000000101110101100111,
24'b000000000101100010110000,
24'b000000000101010100111010,
24'b000000000101000010000010
};
#600;
reall[81] = 0;

pred [81] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 82 False
test_index = 16'd82;
x = {
24'b000000000101100111000111,
24'b000000000101101110010011,
24'b000000000101101101010001,
24'b000000000101011000110000,
24'b000000000101001111100001,
24'b000000000100100110011110,
24'b000000000100011100001101,
24'b000000000100100100011011,
24'b000000000101110101011110,
24'b000000000110000001110010
};
#600;
reall[82] = 0;

pred [82] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 83 False
test_index = 16'd83;
x = {
24'b000000000110000011100000,
24'b000000000110000110100111,
24'b000000000110000110100111,
24'b000000000110000011100000,
24'b000000000110000000011000,
24'b000000000101111101010001,
24'b000000000110001100110101,
24'b000000000110000110100111,
24'b000000000110000101000011,
24'b000000000101111000100110
};
#600;
reall[83] = 0;

pred [83] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 84 False
test_index = 16'd84;
x = {
24'b000000000110101011001110,
24'b000000000110100001001011,
24'b000000000110010001100100,
24'b000000000101111010001001,
24'b000000000101111100010111,
24'b000000000101111110100110,
24'b000000000110000110011010,
24'b000000000101101110111111,
24'b000000000101110110110011,
24'b000000000101111011010000
};
#600;
reall[84] = 0;

pred [84] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 85 True
test_index = 16'd85;
x = {
24'b000000000110011100111111,
24'b000000000110010100100000,
24'b000000000101001111001101,
24'b000000000110111001010010,
24'b000000000111000011001011,
24'b000000000111000110000000,
24'b000000000110110000110010,
24'b000000000110011011100101,
24'b000000000100111001111111,
24'b000000000110101001101110
};
#600;
reall[85] = 1;

pred [85] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 86 False
test_index = 16'd86;
x = {
24'b000000000100011010101111,
24'b000000000100100010011000,
24'b000000000100001100010011,
24'b000000000100010010010000,
24'b000000000100010000100011,
24'b000000000100000010111110,
24'b000000000100010011000110,
24'b000000000100100001100010,
24'b000000000100011111110101,
24'b000000000100000010000111
};
#600;
reall[86] = 0;

pred [86] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 87 False
test_index = 16'd87;
x = {
24'b000000000101101010100010,
24'b000000000101110111010000,
24'b000000000101110000111001,
24'b000000000101111000110110,
24'b000000000101111000110110,
24'b000000000101110000111001,
24'b000000000101100111010110,
24'b000000000101111000110110,
24'b000000000101111101100111,
24'b000000000101110111010000
};
#600;
reall[87] = 0;

pred [87] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 88 True
test_index = 16'd88;
x = {
24'b000000000100111010000010,
24'b000000000001101001101011,
24'b000000000001101001101011,
24'b000000000110010000010111,
24'b000000000100010011010110,
24'b000000000101010111110100,
24'b000000000011110100000101,
24'b000000000011000000000000,
24'b000000000011000001011111,
24'b000000000100111000100011
};
#600;
reall[88] = 1;

pred [88] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 89 False
test_index = 16'd89;
x = {
24'b000000000101100111101000,
24'b000000000101101010011110,
24'b000000000101001111000001,
24'b000000000101100011110110,
24'b000000000101011111000111,
24'b000000000101101100010111,
24'b000000000101000101100011,
24'b000000000101010000111010,
24'b000000000101111111010010,
24'b000000000101110000001001
};
#600;
reall[89] = 0;

pred [89] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 90 False
test_index = 16'd90;
x = {
24'b000000000101110111010000,
24'b000000000101111010011011,
24'b000000000101110010011111,
24'b000000000101100101110000,
24'b000000000101101101101101,
24'b000000000101101101101101,
24'b000000000101110010011111,
24'b000000000101110101101010,
24'b000000000101101000111100,
24'b000000000101101000111100
};
#600;
reall[90] = 0;

pred [90] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 91 False
test_index = 16'd91;
x = {
24'b000000000001011011100000,
24'b000000000010010000101101,
24'b000000000001011110011110,
24'b000000000000111001011101,
24'b000000000001101010011001,
24'b000000000001010110011001,
24'b000000000010000100010111,
24'b000000000010010101110011,
24'b000000000010010010110101,
24'b000000000010001100011100
};
#600;
reall[91] = 0;

pred [91] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 92 False
test_index = 16'd92;
x = {
24'b000000000101101100011100,
24'b000000000101110000111000,
24'b000000000101101100011100,
24'b000000000101110000111000,
24'b000000000101101001011111,
24'b000000000101101000000001,
24'b000000000101110010010110,
24'b000000000101110011110100,
24'b000000000101101000000001,
24'b000000000101100011100110
};
#600;
reall[92] = 0;

pred [92] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 93 False
test_index = 16'd93;
x = {
24'b000000000100110101001110,
24'b000000000100111001000001,
24'b000000000100110010101100,
24'b000000000100101100010110,
24'b000000000100110011111101,
24'b000000000100111111010111,
24'b000000000100110010101100,
24'b000000000100110000001010,
24'b000000000100110000001010,
24'b000000000100110011111101
};
#600;
reall[93] = 0;

pred [93] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 94 False
test_index = 16'd94;
x = {
24'b000000000111011110111001,
24'b000000000111101100001000,
24'b000000000111010010110000,
24'b000000000111100111101110,
24'b000000000111011100101100,
24'b000000000111101110010110,
24'b000000000111100000000000,
24'b000000000111011110111001,
24'b000000000111011011100101,
24'b000000000111001110010110
};
#600;
reall[94] = 0;

pred [94] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 95 True
test_index = 16'd95;
x = {
24'b000000000110110101001111,
24'b000000000010100111100000,
24'b000000000110100010010011,
24'b000000000010101000011101,
24'b000000000010011100001001,
24'b000000000110111010111010,
24'b000000000001011110101000,
24'b000000000001011110101000,
24'b000000000110111001111101,
24'b000000000010101001011001
};
#600;
reall[95] = 1;

pred [95] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 96 False
test_index = 16'd96;
x = {
24'b000000000101101100011100,
24'b000000000101110110110001,
24'b000000000101111100101011,
24'b000000000101111011001101,
24'b000000000101101010111110,
24'b000000000110000001000110,
24'b000000000101110010010110,
24'b000000000101110110110001,
24'b000000000101111111101000,
24'b000000000101111011001101
};
#600;
reall[96] = 0;

pred [96] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 97 True
test_index = 16'd97;
x = {
24'b000000000110110101100111,
24'b000000000100101111010101,
24'b000000000010111100011000,
24'b000000000110101111110100,
24'b000000000100110000010011,
24'b000000000001101011001110,
24'b000000000001100001100100,
24'b000000000110100111000111,
24'b000000000010110101100111,
24'b000000000111001110101110
};
#600;
reall[97] = 1;

pred [97] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 98 False
test_index = 16'd98;
x = {
24'b000000000100011101100000,
24'b000000000100011000101100,
24'b000000000100101111100101,
24'b000000000100010111011111,
24'b000000000100010101000101,
24'b000000000100010011111000,
24'b000000000100100111001001,
24'b000000000100011110101110,
24'b000000000100100011100010,
24'b000000000100011101100000
};
#600;
reall[98] = 0;

pred [98] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
    
// Testcase 99 False
test_index = 16'd99;
x = {
24'b000000000101001001100000,
24'b000000000101001100000010,
24'b000000000101001000001111,
24'b000000000101000101101100,
24'b000000000101000101101100,
24'b000000000101001110100100,
24'b000000000101001000001111,
24'b000000000100111111010111,
24'b000000000101000000101000,
24'b000000000101001000001111
};
#600;
reall[99] = 0;

pred [99] = compare_sign_mag(y1, y2);
reset = 1;
x = 0;
// Wait for global reset to finish
#10;
reset = 0;
        
        // Initialize variables
        sum = 0;
        true = 0;

        for (i = 0; i < max_data; i = i + 1) begin
            if (!(reall[i] === 1'bx || pred[i] === 1'bx)) begin
                $display("testcase: %d, real: %b, pred: %b", i, reall[i], pred[i]);
                sum = sum + 1;
                if (reall[i] == pred[i]) begin
                    true = true + 1;
                end
            end
        end

        if (sum > 0) begin
            $display("accuracy = (%d / %d) = %.3f%%", true, sum, true * 100.0 / sum);
        end else begin
            $display("No valid test cases to calculate accuracy.");
        end

        // Finish simulation
        $finish;
    end

    initial begin
        // // Initialize variables
        // sum = 0;
        // true = 0;

        // for (i = 0; i < 25; i = i + 1) begin
        //     if (!(reall[i] === 1'bx || pred[i] === 1'bx)) begin
        //         $display("testcase: %d, real: %b, pred: %b", i, reall[i], pred[i]);
        //         sum = sum + 1;
        //         if (reall[i] == pred[i]) begin
        //             true = true + 1;
        //         end
        //     end
        // end

        // if (sum > 0) begin
        //     $display("accuracy = %4d / %4d = %4f", true, sum, true * 1.0 / sum);
        // end else begin
        //     $display("No valid test cases to calculate accuracy.");
        // end
    end

endmodule
