`timescale 1ns/1ps
`include "encoder_fixed_point.v"
`include "fixed_point_multiply.v"
`include "fixed_point_add.v"

module tb_encoder_fixed_point;

    // Parameter
    parameter N_input = 9;       // Jumlah input
    parameter M_output = 4;      // Jumlah output
    parameter BITSIZE = 32;      // Ukuran data fixed-point

    // Port untuk modul encoder
    reg [N_input*BITSIZE-1:0] x;         // Flattened input data
    reg [N_input*M_output*BITSIZE-1:0] w; // Flattened weights
    reg [M_output*BITSIZE-1:0] b;       // Flattened biases
    wire [M_output*BITSIZE-1:0] output; // Flattened output

    reg clk;                            // Clock
    reg rst;                            // Reset

    // Instance modul encoder
    encoder_fixed_point #(
        .N_input(N_input),
        .M_output(M_output),
        .BITSIZE(BITSIZE)
    ) encoder_inst (
        .x(x),
        .w(w),
        .b(b),
        .output(output),
        .clk(clk),
        .rst(rst)
    );

    // Clock generation
    always #10 clk = ~clk;

    initial begin
        // Inisialisasi clock dan reset
        clk = 0;
        rst = 1;

        // Reset aktif
        #20;
        rst = 0;

        // Test Case 1
        // Input data: 32-bit fixed-point, flattened
        x = {
            32'b0_01111_000000000000000000000000000, // x[8] = 1.0
            32'b0_01110_100000000000000000000000000, // x[7] = 0.5
            32'b1_01111_000000000000000000000000000, // x[6] = -1.0
            32'b0_01111_000000000000000000000000000, // x[5] = 1.0
            32'b0_01110_100000000000000000000000000, // x[4] = 0.5
            32'b1_01111_000000000000000000000000000, // x[3] = -1.0
            32'b0_01111_000000000000000000000000000, // x[2] = 1.0
            32'b0_01110_100000000000000000000000000, // x[1] = 0.5
            32'b1_01111_000000000000000000000000000  // x[0] = -1.0
        };

        // Bobot: 32-bit fixed-point, flattened
        w = {
            32'b0_01111_000000000000000000000000000, // w[8][3]
            32'b1_01111_000000000000000000000000000, // w[7][3]
            32'b0_01111_000000000000000000000000000, // w[6][3]
            32'b0_01111_000000000000000000000000000, // w[5][3]
            32'b0_01110_100000000000000000000000000, // w[4][3]
            32'b1_01111_000000000000000000000000000, // w[3][3]
            32'b0_01111_000000000000000000000000000, // w[2][3]
            32'b1_01110_100000000000000000000000000, // w[1][3]
            32'b0_01110_100000000000000000000000000, // w[0][3]
            32'b0_01111_000000000000000000000000000, // w[8][2]
            32'b0_01110_100000000000000000000000000, // w[7][2]
            32'b1_01111_000000000000000000000000000, // w[6][2]
            32'b0_01111_000000000000000000000000000, // w[5][2]
            32'b0_01110_100000000000000000000000000, // w[4][2]
            32'b1_01111_000000000000000000000000000, // w[3][2]
            32'b0_01111_000000000000000000000000000, // w[2][2]
            32'b1_01110_100000000000000000000000000, // w[1][2]
            32'b0_01110_100000000000000000000000000, // w[0][2]
            32'b0_01111_000000000000000000000000000, // w[8][1]
            32'b0_01110_100000000000000000000000000, // w[7][1]
            32'b1_01111_000000000000000000000000000, // w[6][1]
            32'b0_01111_000000000000000000000000000, // w[5][1]
            32'b0_01110_100000000000000000000000000, // w[4][1]
            32'b1_01111_000000000000000000000000000, // w[3][1]
            32'b0_01111_000000000000000000000000000, // w[2][1]
            32'b1_01110_100000000000000000000000000, // w[1][1]
            32'b0_01110_100000000000000000000000000, // w[0][1]
            32'b0_01111_000000000000000000000000000, // w[8][0]
            32'b0_01110_100000000000000000000000000, // w[7][0]
            32'b1_01111_000000000000000000000000000, // w[6][0]
            32'b0_01111_000000000000000000000000000, // w[5][0]
            32'b0_01110_100000000000000000000000000, // w[4][0]
            32'b1_01111_000000000000000000000000000, // w[3][0]
            32'b0_01111_000000000000000000000000000, // w[2][0]
            32'b1_01110_100000000000000000000000000, // w[1][0]
            32'b0_01110_100000000000000000000000000  // w[0][0]
        };

        // Biases: 32-bit fixed-point, flattened
        b = {
            32'b1_01111_000000000000000000000000000, // b[3] = -1.0
            32'b0_01111_000000000000000000000000000, // b[2] = 1.0
            32'b0_01110_100000000000000000000000000, // b[1] = 0.5
            32'b0_01111_000000000000000000000000000  // b[0] = 1.0
        };

        // Tunggu beberapa saat untuk hasil
        #100;

        // Stop simulation
        $stop;
    end

    // Monitor output
    initial begin
        $monitor("Time=%0d, Output=%h", $time, output);
    end

endmodule
