`timescale 1ns/1ps
// Basic needs
`include "fixed_point_add.v"
`include "fixed_point_multiply.v"
`include "compare_8float_v2.v"

// Big layer
`include "enc_1.v"
`include "enc_2.v"
// lambda layer
`include "lambda_layer.v"
`include "delay3cc.v"
`include "squareroot.v"
`include "PRNG.v"
// Lanjut big layer
`include "enc_3.v"
`include "enc_4.v"

// enc
`include "enc_control.v"

// Activation function
`include "sigmoid_piped.v"
`include "softplus_8slice_piped.v"

module top_arrhythmia #(parameter BITSIZE = 16) (
    input wire  clk,
    input wire  reset,
    input wire  [BITSIZE*10-1:0]   x,  // Input vector (10 elements)    
    output wire [BITSIZE*2-1:0]    y   // Output vector (2 elements)
);
    // First Layer
    reg signed[BITSIZE*10*6-1:0] w_enc_1;
    reg signed[BITSIZE*6-1:0] b_enc_1;

    initial begin
        w_enc_1 = {
16'b0000000111100111,
16'b0000100010000110,
16'b1000001000101101,
16'b0000000011010110,
16'b0000101010000010,
16'b0000000100101111,
16'b1000001011111110,
16'b1000100001110011,
16'b1000101000100001,
16'b1000010001010011,
16'b0000000001110111,
16'b0000111110000111,
16'b1000000000011001,
16'b0000100111001000,
16'b0000110010111101,
16'b0000000001101001,
16'b0000010111110001,
16'b1001001111000111,
16'b1000000001001101,
16'b1000100010010100,
16'b1000001000100001,
16'b1000000001010010,
16'b0000001101101100,
16'b0000110001000011,
16'b0000000001100101,
16'b0000011100011100,
16'b0000100011010101,
16'b0000000110110110,
16'b0000000000001110,
16'b1001000000000010,
16'b1000000001000110,
16'b1000111111011100,
16'b0000100000111011,
16'b0000000001011011,
16'b0000001010101111,
16'b0000100100110010,
16'b0000001110000100,
16'b0001011011111101,
16'b1001010111101000,
16'b0000001110101011,
16'b0000010011011001,
16'b0000000110001111,
16'b0000000000101010,
16'b1000111110111111,
16'b0000110000000011,
16'b1000000001010101,
16'b0000011011111010,
16'b0000100011100111,
16'b0000000001111000,
16'b0001001001110011,
16'b1000001011010110,
16'b0000000010101100,
16'b0000010110000100,
16'b1000110100111011,
16'b1000000101111101,
16'b1000101001000100,
16'b0000001111110111,
16'b1000000011111110,
16'b0000001000110010,
16'b0000011101110010,
};
b_enc_1 = {
16'b0000000110010111,
16'b1000010011100010,
16'b1000010101101110,
16'b0000000111110111,
16'b0000010011111001,
16'b1000010111010101,
};

    end

endmodule